
module sfilt ( clk, rst, pushin, cmd, q, h, pushout, z );
  input [1:0] cmd;
  input [31:0] q;
  input [31:0] h;
  output [31:0] z;
  input clk, rst, pushin;
  output pushout;
  wire   push1, _pushout_d, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, \C1/DATA1_63 , \C1/DATA1_59 , \C1/DATA1_51 ,
         \C1/DATA1_50 , \C1/DATA1_47 , \C1/DATA1_45 , \C1/DATA1_43 ,
         \C1/DATA1_42 , \C1/DATA1_41 , \C1/DATA1_35 , \C1/DATA1_32 ,
         \C1/DATA1_31 , \C1/DATA1_30 , \C1/DATA1_29 , \C1/DATA1_27 ,
         \C1/DATA1_24 , \C1/DATA1_16 , \C1/DATA1_15 , \C1/DATA1_13 ,
         \C1/DATA1_10 , \C1/DATA1_7 , \C1/DATA1_6 , \C1/DATA1_5 , \C1/DATA1_4 ,
         \C1/DATA1_3 , \C1/DATA1_2 , \C1/DATA1_1 , \C1/DATA1_0 ,
         \DP_OP_14_298_9081/n522 , \DP_OP_14_298_9081/n521 ,
         \DP_OP_14_298_9081/n520 , \DP_OP_14_298_9081/n515 ,
         \DP_OP_14_298_9081/n513 , \DP_OP_14_298_9081/n512 ,
         \DP_OP_14_298_9081/n509 , \DP_OP_14_298_9081/n497 ,
         \DP_OP_14_298_9081/n496 , \DP_OP_14_298_9081/n493 ,
         \DP_OP_14_298_9081/n490 , \DP_OP_14_298_9081/n484 ,
         \DP_OP_14_298_9081/n483 , \DP_OP_14_298_9081/n482 ,
         \DP_OP_14_298_9081/n478 , \DP_OP_14_298_9081/n475 ,
         \DP_OP_14_298_9081/n474 , \DP_OP_14_298_9081/n466 ,
         \DP_OP_14_298_9081/n461 , \DP_OP_14_298_9081/n459 ,
         \DP_OP_14_298_9081/n458 , \DP_OP_14_298_9081/n457 ,
         \DP_OP_14_298_9081/n456 , \DP_OP_14_298_9081/n455 ,
         \DP_OP_14_298_9081/n454 , \DP_OP_14_298_9081/n453 ,
         \DP_OP_14_298_9081/n452 , \DP_OP_14_298_9081/n451 ,
         \DP_OP_14_298_9081/n450 , \DP_OP_14_298_9081/n449 ,
         \DP_OP_14_298_9081/n448 , \DP_OP_14_298_9081/n447 ,
         \DP_OP_14_298_9081/n446 , \DP_OP_14_298_9081/n445 ,
         \DP_OP_14_298_9081/n444 , \DP_OP_14_298_9081/n442 ,
         \DP_OP_14_298_9081/n441 , \DP_OP_14_298_9081/n440 ,
         \DP_OP_14_298_9081/n439 , \DP_OP_14_298_9081/n438 ,
         \DP_OP_14_298_9081/n437 , \DP_OP_14_298_9081/n436 ,
         \DP_OP_14_298_9081/n435 , \DP_OP_14_298_9081/n434 ,
         \DP_OP_14_298_9081/n433 , \DP_OP_14_298_9081/n432 ,
         \DP_OP_14_298_9081/n431 , \DP_OP_14_298_9081/n430 ,
         \DP_OP_14_298_9081/n429 , \DP_OP_14_298_9081/n428 ,
         \DP_OP_14_298_9081/n427 , \DP_OP_14_298_9081/n426 ,
         \DP_OP_14_298_9081/n425 , \DP_OP_14_298_9081/n424 ,
         \DP_OP_14_298_9081/n422 , \DP_OP_14_298_9081/n421 ,
         \DP_OP_14_298_9081/n420 , \DP_OP_14_298_9081/n419 ,
         \DP_OP_14_298_9081/n418 , \DP_OP_14_298_9081/n417 ,
         \DP_OP_14_298_9081/n416 , \DP_OP_14_298_9081/n415 ,
         \DP_OP_14_298_9081/n414 , \DP_OP_14_298_9081/n410 ,
         \DP_OP_14_298_9081/n409 , \DP_OP_14_298_9081/n408 ,
         \DP_OP_14_298_9081/n407 , \DP_OP_14_298_9081/n406 ,
         \DP_OP_14_298_9081/n405 , \DP_OP_14_298_9081/n404 ,
         \DP_OP_14_298_9081/n403 , \DP_OP_14_298_9081/n402 ,
         \DP_OP_14_298_9081/n401 , \DP_OP_14_298_9081/n399 ,
         \DP_OP_14_298_9081/n398 , \DP_OP_14_298_9081/n397 ,
         \DP_OP_14_298_9081/n396 , \DP_OP_14_298_9081/n395 ,
         \DP_OP_14_298_9081/n394 , \DP_OP_14_298_9081/n393 ,
         \DP_OP_14_298_9081/n392 , \DP_OP_14_298_9081/n390 ,
         \DP_OP_14_298_9081/n389 , \DP_OP_14_298_9081/n388 ,
         \DP_OP_14_298_9081/n387 , \DP_OP_14_298_9081/n386 ,
         \DP_OP_14_298_9081/n385 , \DP_OP_14_298_9081/n384 ,
         \DP_OP_14_298_9081/n383 , \DP_OP_14_298_9081/n381 ,
         \DP_OP_14_298_9081/n380 , \DP_OP_14_298_9081/n379 ,
         \DP_OP_14_298_9081/n375 , \DP_OP_14_298_9081/n374 ,
         \DP_OP_14_298_9081/n373 , \DP_OP_14_298_9081/n372 ,
         \DP_OP_14_298_9081/n371 , \DP_OP_14_298_9081/n370 ,
         \DP_OP_14_298_9081/n369 , \DP_OP_14_298_9081/n367 ,
         \DP_OP_14_298_9081/n366 , \DP_OP_14_298_9081/n365 ,
         \DP_OP_14_298_9081/n364 , \DP_OP_14_298_9081/n363 ,
         \DP_OP_14_298_9081/n362 , \DP_OP_14_298_9081/n361 ,
         \DP_OP_14_298_9081/n360 , \DP_OP_14_298_9081/n359 ,
         \DP_OP_14_298_9081/n358 , \DP_OP_14_298_9081/n356 ,
         \DP_OP_14_298_9081/n355 , \DP_OP_14_298_9081/n354 ,
         \DP_OP_14_298_9081/n353 , \DP_OP_14_298_9081/n352 ,
         \DP_OP_14_298_9081/n351 , \DP_OP_14_298_9081/n350 ,
         \DP_OP_14_298_9081/n348 , \DP_OP_14_298_9081/n347 ,
         \DP_OP_14_298_9081/n346 , \DP_OP_14_298_9081/n345 ,
         \DP_OP_14_298_9081/n344 , \DP_OP_14_298_9081/n343 ,
         \DP_OP_14_298_9081/n342 , \DP_OP_14_298_9081/n341 ,
         \DP_OP_14_298_9081/n340 , \DP_OP_14_298_9081/n339 ,
         \DP_OP_14_298_9081/n338 , \DP_OP_14_298_9081/n337 ,
         \DP_OP_14_298_9081/n336 , \DP_OP_14_298_9081/n335 ,
         \DP_OP_14_298_9081/n333 , \DP_OP_14_298_9081/n332 ,
         \DP_OP_14_298_9081/n331 , \DP_OP_14_298_9081/n330 ,
         \DP_OP_14_298_9081/n329 , \DP_OP_14_298_9081/n328 ,
         \DP_OP_14_298_9081/n327 , \DP_OP_14_298_9081/n325 ,
         \DP_OP_14_298_9081/n324 , \DP_OP_14_298_9081/n323 ,
         \DP_OP_14_298_9081/n322 , \DP_OP_14_298_9081/n321 ,
         \DP_OP_14_298_9081/n320 , \DP_OP_14_298_9081/n319 ,
         \DP_OP_14_298_9081/n318 , \DP_OP_14_298_9081/n317 ,
         \DP_OP_14_298_9081/n316 , \DP_OP_14_298_9081/n315 ,
         \DP_OP_14_298_9081/n314 , \DP_OP_14_298_9081/n313 ,
         \DP_OP_14_298_9081/n312 , \DP_OP_14_298_9081/n310 ,
         \DP_OP_14_298_9081/n309 , \DP_OP_14_298_9081/n308 ,
         \DP_OP_14_298_9081/n307 , \DP_OP_14_298_9081/n306 ,
         \DP_OP_14_298_9081/n305 , \DP_OP_14_298_9081/n304 ,
         \DP_OP_14_298_9081/n303 , \DP_OP_14_298_9081/n301 ,
         \DP_OP_14_298_9081/n300 , \DP_OP_14_298_9081/n299 ,
         \DP_OP_14_298_9081/n298 , \DP_OP_14_298_9081/n297 ,
         \DP_OP_14_298_9081/n296 , \DP_OP_14_298_9081/n295 ,
         \DP_OP_14_298_9081/n294 , \DP_OP_14_298_9081/n293 ,
         \DP_OP_14_298_9081/n292 , \DP_OP_14_298_9081/n290 ,
         \DP_OP_14_298_9081/n289 , \DP_OP_14_298_9081/n288 ,
         \DP_OP_14_298_9081/n286 , \DP_OP_14_298_9081/n285 ,
         \DP_OP_14_298_9081/n284 , \DP_OP_14_298_9081/n283 ,
         \DP_OP_14_298_9081/n282 , \DP_OP_14_298_9081/n281 ,
         \DP_OP_14_298_9081/n280 , \DP_OP_14_298_9081/n279 ,
         \DP_OP_14_298_9081/n278 , \DP_OP_14_298_9081/n277 ,
         \DP_OP_14_298_9081/n276 , \DP_OP_14_298_9081/n275 ,
         \DP_OP_14_298_9081/n270 , \DP_OP_14_298_9081/n269 ,
         \DP_OP_14_298_9081/n268 , \DP_OP_14_298_9081/n267 ,
         \DP_OP_14_298_9081/n266 , \DP_OP_14_298_9081/n265 ,
         \DP_OP_14_298_9081/n264 , \DP_OP_14_298_9081/n262 ,
         \DP_OP_14_298_9081/n261 , \DP_OP_14_298_9081/n260 ,
         \DP_OP_14_298_9081/n259 , \DP_OP_14_298_9081/n258 ,
         \DP_OP_14_298_9081/n257 , \DP_OP_14_298_9081/n256 ,
         \DP_OP_14_298_9081/n255 , \DP_OP_14_298_9081/n254 ,
         \DP_OP_14_298_9081/n253 , \DP_OP_14_298_9081/n252 ,
         \DP_OP_14_298_9081/n250 , \DP_OP_14_298_9081/n249 ,
         \DP_OP_14_298_9081/n248 , \DP_OP_14_298_9081/n247 ,
         \DP_OP_14_298_9081/n246 , \DP_OP_14_298_9081/n245 ,
         \DP_OP_14_298_9081/n242 , \DP_OP_14_298_9081/n241 ,
         \DP_OP_14_298_9081/n240 , \DP_OP_14_298_9081/n239 ,
         \DP_OP_14_298_9081/n238 , \DP_OP_14_298_9081/n237 ,
         \DP_OP_14_298_9081/n236 , \DP_OP_14_298_9081/n235 ,
         \DP_OP_14_298_9081/n234 , \DP_OP_14_298_9081/n233 ,
         \DP_OP_14_298_9081/n232 , \DP_OP_14_298_9081/n231 ,
         \DP_OP_14_298_9081/n230 , \DP_OP_14_298_9081/n229 ,
         \DP_OP_14_298_9081/n228 , \DP_OP_14_298_9081/n227 ,
         \DP_OP_14_298_9081/n226 , \DP_OP_14_298_9081/n225 ,
         \DP_OP_14_298_9081/n224 , \DP_OP_14_298_9081/n223 ,
         \DP_OP_14_298_9081/n222 , \DP_OP_14_298_9081/n221 ,
         \DP_OP_14_298_9081/n220 , \DP_OP_14_298_9081/n219 ,
         \DP_OP_14_298_9081/n218 , \DP_OP_14_298_9081/n217 ,
         \DP_OP_14_298_9081/n216 , \DP_OP_14_298_9081/n215 ,
         \DP_OP_14_298_9081/n214 , \DP_OP_14_298_9081/n213 ,
         \DP_OP_14_298_9081/n212 , \DP_OP_14_298_9081/n211 ,
         \DP_OP_14_298_9081/n210 , \DP_OP_14_298_9081/n209 ,
         \DP_OP_14_298_9081/n208 , \DP_OP_14_298_9081/n206 ,
         \DP_OP_14_298_9081/n205 , \DP_OP_14_298_9081/n204 ,
         \DP_OP_14_298_9081/n203 , \DP_OP_14_298_9081/n202 ,
         \DP_OP_14_298_9081/n201 , \DP_OP_14_298_9081/n200 ,
         \DP_OP_14_298_9081/n199 , \DP_OP_14_298_9081/n198 ,
         \DP_OP_14_298_9081/n197 , \DP_OP_14_298_9081/n196 ,
         \DP_OP_14_298_9081/n195 , \DP_OP_14_298_9081/n194 ,
         \DP_OP_14_298_9081/n193 , \DP_OP_14_298_9081/n192 ,
         \DP_OP_14_298_9081/n191 , \DP_OP_14_298_9081/n190 ,
         \DP_OP_14_298_9081/n189 , \DP_OP_14_298_9081/n188 ,
         \DP_OP_14_298_9081/n187 , \DP_OP_14_298_9081/n184 ,
         \DP_OP_14_298_9081/n183 , \DP_OP_14_298_9081/n182 ,
         \DP_OP_14_298_9081/n181 , \DP_OP_14_298_9081/n180 ,
         \DP_OP_14_298_9081/n178 , \DP_OP_14_298_9081/n177 ,
         \DP_OP_14_298_9081/n176 , \DP_OP_14_298_9081/n175 ,
         \DP_OP_14_298_9081/n174 , \DP_OP_14_298_9081/n173 ,
         \DP_OP_14_298_9081/n172 , \DP_OP_14_298_9081/n171 ,
         \DP_OP_14_298_9081/n170 , \DP_OP_14_298_9081/n169 ,
         \DP_OP_14_298_9081/n168 , \DP_OP_14_298_9081/n167 ,
         \DP_OP_14_298_9081/n166 , \DP_OP_14_298_9081/n165 ,
         \DP_OP_14_298_9081/n164 , \DP_OP_14_298_9081/n163 ,
         \DP_OP_14_298_9081/n160 , \DP_OP_14_298_9081/n159 ,
         \DP_OP_14_298_9081/n158 , \DP_OP_14_298_9081/n157 ,
         \DP_OP_14_298_9081/n156 , \DP_OP_14_298_9081/n155 ,
         \DP_OP_14_298_9081/n154 , \DP_OP_14_298_9081/n153 ,
         \DP_OP_14_298_9081/n152 , \DP_OP_14_298_9081/n150 ,
         \DP_OP_14_298_9081/n149 , \DP_OP_14_298_9081/n148 ,
         \DP_OP_14_298_9081/n145 , \DP_OP_14_298_9081/n144 ,
         \DP_OP_14_298_9081/n143 , \DP_OP_14_298_9081/n142 ,
         \DP_OP_14_298_9081/n141 , \DP_OP_14_298_9081/n140 ,
         \DP_OP_14_298_9081/n139 , \DP_OP_14_298_9081/n138 ,
         \DP_OP_14_298_9081/n136 , \DP_OP_14_298_9081/n135 ,
         \DP_OP_14_298_9081/n134 , \DP_OP_14_298_9081/n133 ,
         \DP_OP_14_298_9081/n132 , \DP_OP_14_298_9081/n131 ,
         \DP_OP_14_298_9081/n130 , \DP_OP_14_298_9081/n129 ,
         \DP_OP_14_298_9081/n128 , \DP_OP_14_298_9081/n127 ,
         \DP_OP_14_298_9081/n126 , \DP_OP_14_298_9081/n125 ,
         \DP_OP_14_298_9081/n124 , \DP_OP_14_298_9081/n123 ,
         \DP_OP_14_298_9081/n122 , \DP_OP_14_298_9081/n120 ,
         \DP_OP_14_298_9081/n119 , \DP_OP_14_298_9081/n118 ,
         \DP_OP_14_298_9081/n115 , \DP_OP_14_298_9081/n114 ,
         \DP_OP_14_298_9081/n113 , \DP_OP_14_298_9081/n112 ,
         \DP_OP_14_298_9081/n111 , \DP_OP_14_298_9081/n110 ,
         \DP_OP_14_298_9081/n109 , \DP_OP_14_298_9081/n108 ,
         \DP_OP_14_298_9081/n107 , \DP_OP_14_298_9081/n106 ,
         \DP_OP_14_298_9081/n105 , \DP_OP_14_298_9081/n104 ,
         \DP_OP_14_298_9081/n103 , \DP_OP_14_298_9081/n102 ,
         \DP_OP_14_298_9081/n101 , \DP_OP_14_298_9081/n100 ,
         \DP_OP_14_298_9081/n99 , \DP_OP_14_298_9081/n98 ,
         \DP_OP_14_298_9081/n97 , \DP_OP_14_298_9081/n96 ,
         \DP_OP_14_298_9081/n95 , \DP_OP_14_298_9081/n94 ,
         \DP_OP_14_298_9081/n91 , \DP_OP_14_298_9081/n90 ,
         \DP_OP_14_298_9081/n89 , \DP_OP_14_298_9081/n88 ,
         \DP_OP_14_298_9081/n86 , \DP_OP_14_298_9081/n84 ,
         \DP_OP_14_298_9081/n82 , \DP_OP_14_298_9081/n81 ,
         \DP_OP_14_298_9081/n80 , \DP_OP_14_298_9081/n79 ,
         \DP_OP_14_298_9081/n78 , \DP_OP_14_298_9081/n77 ,
         \DP_OP_14_298_9081/n76 , \DP_OP_14_298_9081/n75 ,
         \DP_OP_14_298_9081/n74 , \DP_OP_14_298_9081/n73 ,
         \DP_OP_14_298_9081/n72 , \DP_OP_14_298_9081/n71 ,
         \DP_OP_14_298_9081/n70 , \DP_OP_14_298_9081/n67 ,
         \DP_OP_14_298_9081/n65 , \DP_OP_14_298_9081/n64 ,
         \DP_OP_14_298_9081/n63 , \DP_OP_14_298_9081/n61 ,
         \DP_OP_14_298_9081/n58 , \DP_OP_14_298_9081/n55 ,
         \DP_OP_14_298_9081/n52 , \DP_OP_14_298_9081/n39 ,
         \DP_OP_14_298_9081/n36 , \DP_OP_14_298_9081/n33 ,
         \DP_OP_14_298_9081/n27 , \DP_OP_14_298_9081/n26 ,
         \DP_OP_14_298_9081/n25 , \DP_OP_14_298_9081/n21 ,
         \DP_OP_14_298_9081/n18 , \DP_OP_14_298_9081/n17 ,
         \DP_OP_14_298_9081/n9 , \DP_OP_14_298_9081/n5 ,
         \DP_OP_14_298_9081/n4 , \DP_OP_14_298_9081/n3 ,
         \DP_OP_14_298_9081/n2 , \DP_OP_14_298_9081/n1 ,
         \DP_OP_14_298_9081/n487 , \DP_OP_14_298_9081/n30 , \C1/DATA1_38 ,
         \DP_OP_14_298_9081/n468 , \DP_OP_14_298_9081/n121 ,
         \DP_OP_14_298_9081/n11 , \C1/DATA1_57 , \DP_OP_14_298_9081/n473 ,
         \DP_OP_14_298_9081/n16 , \C1/DATA1_52 , \DP_OP_14_298_9081/n470 ,
         \DP_OP_14_298_9081/n137 , \DP_OP_14_298_9081/n13 , \C1/DATA1_55 ,
         \DP_OP_14_298_9081/n6 , \DP_OP_14_298_9081/n463 , \C1/DATA1_62 ,
         \DP_OP_14_298_9081/n485 , \DP_OP_14_298_9081/n28 , \C1/DATA1_40 ,
         \C1/DATA1_11 , \DP_OP_14_298_9081/n481 , \DP_OP_14_298_9081/n24 ,
         \C1/DATA1_44 , \DP_OP_14_298_9081/n467 , \DP_OP_14_298_9081/n10 ,
         \C1/DATA1_58 , \DP_OP_14_298_9081/n472 , \DP_OP_14_298_9081/n151 ,
         \DP_OP_14_298_9081/n15 , \C1/DATA1_53 , \DP_OP_14_298_9081/n8 ,
         \C1/DATA1_60 , \DP_OP_14_298_9081/n477 , \DP_OP_14_298_9081/n20 ,
         \C1/DATA1_48 , \DP_OP_14_298_9081/n476 , \DP_OP_14_298_9081/n19 ,
         \DP_OP_14_298_9081/n179 , \C1/DATA1_49 , \C1/DATA1_25 ,
         \DP_OP_14_298_9081/n488 , \DP_OP_14_298_9081/n31 ,
         \DP_OP_14_298_9081/n263 , \C1/DATA1_37 , \DP_OP_14_298_9081/n492 ,
         \DP_OP_14_298_9081/n35 , \DP_OP_14_298_9081/n287 , \C1/DATA1_33 ,
         \C1/DATA1_20 , \DP_OP_14_298_9081/n469 , \DP_OP_14_298_9081/n12 ,
         \C1/DATA1_56 , \DP_OP_14_298_9081/n87 , \DP_OP_14_298_9081/n7 ,
         \C1/DATA1_61 , \DP_OP_14_298_9081/n471 , \DP_OP_14_298_9081/n14 ,
         \C1/DATA1_54 , n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933;
  wire   [63:0] acc;
  wire   [63:0] acc_a;
  wire   [1:0] cmd1;
  wire   [1:0] cmd2;
  wire   [31:0] q0;
  wire   [31:0] h0;
  wire   [6:0] ho_2;
  wire   [1:0] cmd0;
  wire   [6:0] h0_d_a;
  tri   clk;
  tri   [31:0] q0_d;
  tri   [31:0] h0_d;
  tri   [63:0] out;
  tri   n1934;

  DW02_mult_3_stage a1 ( .A(q0_d), .B(h0_d), .CLK(clk), .TC(1'b1), .PRODUCT(
        out) );
  CFD2QX1 \cmd2_reg[1]  ( .D(n417), .CP(clk), .CD(n199), .Q(cmd2[1]) );
  CFD2QX1 \cmd2_reg[0]  ( .D(n600), .CP(clk), .CD(n199), .Q(cmd2[0]) );
  CFD2QX1 \acc_a_reg[59]  ( .D(n599), .CP(clk), .CD(n199), .Q(acc_a[59]) );
  CFD2QX1 \acc_a_reg[58]  ( .D(n598), .CP(clk), .CD(n199), .Q(acc_a[58]) );
  CFD2QX1 \acc_a_reg[57]  ( .D(n597), .CP(clk), .CD(n199), .Q(acc_a[57]) );
  CFD2QX1 \acc_a_reg[55]  ( .D(n596), .CP(clk), .CD(n199), .Q(acc_a[55]) );
  CFD2QX1 \acc_a_reg[54]  ( .D(n595), .CP(clk), .CD(n199), .Q(acc_a[54]) );
  CFD2QX1 \acc_a_reg[53]  ( .D(n594), .CP(clk), .CD(n199), .Q(acc_a[53]) );
  CFD2QX1 \acc_a_reg[51]  ( .D(n593), .CP(clk), .CD(n199), .Q(acc_a[51]) );
  CFD2QX1 \acc_a_reg[50]  ( .D(n592), .CP(clk), .CD(n199), .Q(acc_a[50]) );
  CFD2QX1 \acc_a_reg[49]  ( .D(n591), .CP(clk), .CD(n199), .Q(acc_a[49]) );
  CFD2QX1 \acc_a_reg[48]  ( .D(n590), .CP(clk), .CD(n199), .Q(acc_a[48]) );
  CFD2QX1 \acc_a_reg[47]  ( .D(n589), .CP(clk), .CD(n199), .Q(acc_a[47]) );
  CFD2QX1 \acc_a_reg[46]  ( .D(n588), .CP(clk), .CD(n199), .Q(acc_a[46]) );
  CFD2QX1 \acc_a_reg[45]  ( .D(n587), .CP(clk), .CD(n199), .Q(acc_a[45]) );
  CFD2QX1 \acc_a_reg[44]  ( .D(n586), .CP(clk), .CD(n199), .Q(acc_a[44]) );
  CFD2QX1 \acc_a_reg[43]  ( .D(n585), .CP(clk), .CD(n199), .Q(acc_a[43]) );
  CFD2QX1 \acc_a_reg[42]  ( .D(n584), .CP(clk), .CD(n199), .Q(acc_a[42]) );
  CFD2QX1 \acc_a_reg[41]  ( .D(n583), .CP(clk), .CD(n199), .Q(acc_a[41]) );
  CFD2QX1 \acc_a_reg[40]  ( .D(n582), .CP(clk), .CD(n199), .Q(acc_a[40]) );
  CFD2QX1 \acc_a_reg[39]  ( .D(n581), .CP(clk), .CD(n199), .Q(acc_a[39]) );
  CFD2QX1 \acc_a_reg[38]  ( .D(n580), .CP(clk), .CD(n199), .Q(acc_a[38]) );
  CFD2QX1 \acc_a_reg[37]  ( .D(n579), .CP(clk), .CD(n199), .Q(acc_a[37]) );
  CFD2QX1 \acc_a_reg[36]  ( .D(n578), .CP(clk), .CD(n199), .Q(acc_a[36]) );
  CFD2QX1 \acc_a_reg[35]  ( .D(n577), .CP(clk), .CD(n199), .Q(acc_a[35]) );
  CFD2QX1 \acc_a_reg[34]  ( .D(n576), .CP(clk), .CD(n199), .Q(acc_a[34]) );
  CFD2QX1 \acc_a_reg[33]  ( .D(n575), .CP(clk), .CD(n199), .Q(acc_a[33]) );
  CFD2QX1 \acc_a_reg[32]  ( .D(n574), .CP(clk), .CD(n199), .Q(acc_a[32]) );
  CFD2QX1 \acc_a_reg[31]  ( .D(n573), .CP(clk), .CD(n199), .Q(acc_a[31]) );
  CFD2QX1 \acc_a_reg[30]  ( .D(n572), .CP(clk), .CD(n199), .Q(acc_a[30]) );
  CFD2QX1 \acc_a_reg[29]  ( .D(n571), .CP(clk), .CD(n199), .Q(acc_a[29]) );
  CFD2QX1 \acc_a_reg[28]  ( .D(n570), .CP(clk), .CD(n199), .Q(acc_a[28]) );
  CFD2QX1 \acc_a_reg[27]  ( .D(n569), .CP(clk), .CD(n199), .Q(acc_a[27]) );
  CFD2QX1 \acc_a_reg[26]  ( .D(n568), .CP(clk), .CD(n199), .Q(acc_a[26]) );
  CFD2QX1 \acc_a_reg[25]  ( .D(n567), .CP(clk), .CD(n199), .Q(acc_a[25]) );
  CFD2QX1 \acc_a_reg[24]  ( .D(n566), .CP(clk), .CD(n199), .Q(acc_a[24]) );
  CFD2QX1 \acc_a_reg[22]  ( .D(n565), .CP(clk), .CD(n199), .Q(acc_a[22]) );
  CFD2QX1 \acc_a_reg[21]  ( .D(n564), .CP(clk), .CD(n199), .Q(acc_a[21]) );
  CFD2QX1 \acc_a_reg[20]  ( .D(n563), .CP(clk), .CD(n199), .Q(acc_a[20]) );
  CFD2QX1 \acc_a_reg[19]  ( .D(n562), .CP(clk), .CD(n199), .Q(acc_a[19]) );
  CFD2QX1 \acc_a_reg[18]  ( .D(n561), .CP(clk), .CD(n199), .Q(acc_a[18]) );
  CFD2QX1 \acc_a_reg[17]  ( .D(n560), .CP(clk), .CD(n199), .Q(acc_a[17]) );
  CFD2QX1 \acc_a_reg[16]  ( .D(n559), .CP(clk), .CD(n199), .Q(acc_a[16]) );
  CFD2QX1 \acc_a_reg[15]  ( .D(n558), .CP(clk), .CD(n199), .Q(acc_a[15]) );
  CFD2QX1 \acc_a_reg[14]  ( .D(n249), .CP(clk), .CD(n199), .Q(acc_a[14]) );
  CFD2QX1 \acc_a_reg[13]  ( .D(n248), .CP(clk), .CD(n199), .Q(acc_a[13]) );
  CFD2QX1 \acc_a_reg[12]  ( .D(n247), .CP(clk), .CD(n199), .Q(acc_a[12]) );
  CFD2QX1 \acc_a_reg[11]  ( .D(n246), .CP(clk), .CD(n199), .Q(acc_a[11]) );
  CFD2QX1 \acc_a_reg[10]  ( .D(n245), .CP(clk), .CD(n199), .Q(acc_a[10]) );
  CFD2QX1 \acc_a_reg[9]  ( .D(n244), .CP(clk), .CD(n199), .Q(acc_a[9]) );
  CFD2QX1 \acc_a_reg[8]  ( .D(n243), .CP(clk), .CD(n199), .Q(acc_a[8]) );
  CFD2QX1 \acc_a_reg[7]  ( .D(n242), .CP(clk), .CD(n199), .Q(acc_a[7]) );
  CFD2QX1 \acc_a_reg[6]  ( .D(n241), .CP(clk), .CD(n199), .Q(acc_a[6]) );
  CFD2QX1 \acc_a_reg[5]  ( .D(n240), .CP(clk), .CD(n199), .Q(acc_a[5]) );
  CFD2QX1 \acc_a_reg[4]  ( .D(n239), .CP(clk), .CD(n199), .Q(acc_a[4]) );
  CFD2QX1 \acc_a_reg[3]  ( .D(n238), .CP(clk), .CD(n199), .Q(acc_a[3]) );
  CFD2QX1 \acc_a_reg[2]  ( .D(n237), .CP(clk), .CD(n199), .Q(acc_a[2]) );
  CFD2QX1 \acc_a_reg[1]  ( .D(n236), .CP(clk), .CD(n199), .Q(acc_a[1]) );
  CFD2QX1 \acc_a_reg[0]  ( .D(n235), .CP(clk), .CD(n199), .Q(acc_a[0]) );
  CFD2QX1 \acc_reg[0]  ( .D(n689), .CP(clk), .CD(n199), .Q(acc[0]) );
  CFD2QX1 \acc_reg[1]  ( .D(n195), .CP(clk), .CD(n199), .Q(acc[1]) );
  CFD2QX1 \acc_reg[4]  ( .D(n192), .CP(clk), .CD(n199), .Q(acc[4]) );
  CFD2QX1 \acc_reg[5]  ( .D(n191), .CP(clk), .CD(n199), .Q(acc[5]) );
  CFD2QX1 \acc_reg[6]  ( .D(n190), .CP(clk), .CD(n199), .Q(acc[6]) );
  CFD2QX1 \acc_reg[7]  ( .D(n189), .CP(clk), .CD(n199), .Q(acc[7]) );
  CFD2QX1 \acc_reg[10]  ( .D(n186), .CP(clk), .CD(n199), .Q(acc[10]) );
  CFD2QX1 \acc_reg[26]  ( .D(n170), .CP(clk), .CD(n199), .Q(acc[26]) );
  CFD2QX1 \acc_reg[27]  ( .D(n169), .CP(clk), .CD(n199), .Q(acc[27]) );
  CFD2QX1 \acc_reg[28]  ( .D(n168), .CP(clk), .CD(n199), .Q(acc[28]) );
  CFD2QX1 \acc_reg[29]  ( .D(n167), .CP(clk), .CD(n199), .Q(acc[29]) );
  CFD2QX1 \acc_reg[30]  ( .D(n166), .CP(clk), .CD(n199), .Q(acc[30]) );
  CFD2QX1 \acc_reg[34]  ( .D(n162), .CP(clk), .CD(n199), .Q(acc[34]) );
  CFD2QX1 \acc_reg[39]  ( .D(n157), .CP(clk), .CD(n199), .Q(acc[39]) );
  CFD2QX1 \acc_reg[46]  ( .D(n150), .CP(clk), .CD(n199), .Q(acc[46]) );
  CFD2QX1 \acc_reg[63]  ( .D(n133), .CP(clk), .CD(n199), .Q(acc[63]) );
  CFD2QX1 \ho_2_reg[6]  ( .D(n553), .CP(clk), .CD(n199), .Q(ho_2[6]) );
  CFD2QX1 \ho_2_reg[5]  ( .D(n552), .CP(clk), .CD(n199), .Q(ho_2[5]) );
  CAOR2X1 U361 ( .A(pushin), .B(q[3]), .C(n1431), .D(q0[3]), .Z(q0_d[3]) );
  CAOR2X1 U362 ( .A(pushin), .B(q[2]), .C(n1432), .D(q0[2]), .Z(q0_d[2]) );
  CAOR2X1 U363 ( .A(pushin), .B(q[1]), .C(n1432), .D(q0[1]), .Z(q0_d[1]) );
  CFD2QX2 \acc_reg[12]  ( .D(n184), .CP(clk), .CD(n199), .Q(acc[12]) );
  CFD2QX2 \ho_2_reg[3]  ( .D(n601), .CP(clk), .CD(n199), .Q(ho_2[3]) );
  CFD2QXL _pushout_reg ( .D(n602), .CP(clk), .CD(n199), .Q(pushout) );
  CFD2QXL \dout_reg[12]  ( .D(n222), .CP(clk), .CD(n199), .Q(z[12]) );
  CFD2QXL \q0_reg[0]  ( .D(n703), .CP(clk), .CD(n199), .Q(q0[0]) );
  CFD2QXL \h0_reg[7]  ( .D(n704), .CP(clk), .CD(n199), .Q(h0[7]) );
  CFD2QXL \h0_reg[8]  ( .D(n705), .CP(clk), .CD(n199), .Q(h0[8]) );
  CFD2QXL \h0_reg[9]  ( .D(n706), .CP(clk), .CD(n199), .Q(h0[9]) );
  CFD2QXL \h0_reg[10]  ( .D(n707), .CP(clk), .CD(n199), .Q(h0[10]) );
  CFD2QXL \h0_reg[11]  ( .D(n708), .CP(clk), .CD(n199), .Q(h0[11]) );
  CFD2QXL \h0_reg[12]  ( .D(n709), .CP(clk), .CD(n199), .Q(h0[12]) );
  CFD2QXL \h0_reg[13]  ( .D(n710), .CP(clk), .CD(n199), .Q(h0[13]) );
  CFD2QXL \h0_reg[14]  ( .D(n711), .CP(clk), .CD(n199), .Q(h0[14]) );
  CFD2QXL \h0_reg[15]  ( .D(n712), .CP(clk), .CD(n199), .Q(h0[15]) );
  CFD2QXL \h0_reg[16]  ( .D(n713), .CP(clk), .CD(n199), .Q(h0[16]) );
  CFD2QXL \h0_reg[17]  ( .D(n714), .CP(clk), .CD(n199), .Q(h0[17]) );
  CFD2QXL \h0_reg[18]  ( .D(n715), .CP(clk), .CD(n199), .Q(h0[18]) );
  CFD2QXL \h0_reg[19]  ( .D(n716), .CP(clk), .CD(n199), .Q(h0[19]) );
  CFD2QXL \h0_reg[20]  ( .D(n717), .CP(clk), .CD(n199), .Q(h0[20]) );
  CFD2QXL \h0_reg[21]  ( .D(n718), .CP(clk), .CD(n199), .Q(h0[21]) );
  CFD2QXL \h0_reg[22]  ( .D(n719), .CP(clk), .CD(n199), .Q(h0[22]) );
  CFD2QXL \h0_reg[23]  ( .D(n720), .CP(clk), .CD(n199), .Q(h0[23]) );
  CFD2QXL \h0_reg[24]  ( .D(n721), .CP(clk), .CD(n199), .Q(h0[24]) );
  CFD2QXL \h0_reg[25]  ( .D(n722), .CP(clk), .CD(n199), .Q(h0[25]) );
  CFD2QXL \h0_reg[26]  ( .D(n723), .CP(clk), .CD(n199), .Q(h0[26]) );
  CFD2QXL \h0_reg[27]  ( .D(n724), .CP(clk), .CD(n199), .Q(h0[27]) );
  CFD2QXL \h0_reg[28]  ( .D(n725), .CP(clk), .CD(n199), .Q(h0[28]) );
  CFD2QXL \h0_reg[29]  ( .D(n726), .CP(clk), .CD(n199), .Q(h0[29]) );
  CFD2QXL \h0_reg[30]  ( .D(n727), .CP(clk), .CD(n199), .Q(h0[30]) );
  CFD2QXL \h0_reg[31]  ( .D(n728), .CP(clk), .CD(n199), .Q(h0[31]) );
  CFD2QXL \q0_reg[1]  ( .D(n729), .CP(clk), .CD(n199), .Q(q0[1]) );
  CFD2QXL \q0_reg[2]  ( .D(n730), .CP(clk), .CD(n199), .Q(q0[2]) );
  CFD2QXL \q0_reg[3]  ( .D(n731), .CP(clk), .CD(n199), .Q(q0[3]) );
  CFD2QXL \q0_reg[4]  ( .D(n732), .CP(clk), .CD(n199), .Q(q0[4]) );
  CFD2QXL \q0_reg[5]  ( .D(n733), .CP(clk), .CD(n199), .Q(q0[5]) );
  CFD2QXL \q0_reg[6]  ( .D(n734), .CP(clk), .CD(n199), .Q(q0[6]) );
  CFD2QXL \q0_reg[7]  ( .D(n735), .CP(clk), .CD(n199), .Q(q0[7]) );
  CFD2QXL \q0_reg[8]  ( .D(n736), .CP(clk), .CD(n199), .Q(q0[8]) );
  CFD2QXL \q0_reg[9]  ( .D(n737), .CP(clk), .CD(n199), .Q(q0[9]) );
  CFD2QXL \q0_reg[10]  ( .D(n738), .CP(clk), .CD(n199), .Q(q0[10]) );
  CFD2QXL \q0_reg[11]  ( .D(n739), .CP(clk), .CD(n199), .Q(q0[11]) );
  CFD2QXL \q0_reg[12]  ( .D(n740), .CP(clk), .CD(n199), .Q(q0[12]) );
  CFD2QXL \q0_reg[13]  ( .D(n741), .CP(clk), .CD(n199), .Q(q0[13]) );
  CFD2QXL \q0_reg[14]  ( .D(n742), .CP(clk), .CD(n199), .Q(q0[14]) );
  CFD2QXL \q0_reg[15]  ( .D(n743), .CP(clk), .CD(n199), .Q(q0[15]) );
  CFD2QXL \q0_reg[16]  ( .D(n744), .CP(clk), .CD(n199), .Q(q0[16]) );
  CFD2QXL \q0_reg[17]  ( .D(n745), .CP(clk), .CD(n199), .Q(q0[17]) );
  CFD2QXL \q0_reg[18]  ( .D(n746), .CP(clk), .CD(n199), .Q(q0[18]) );
  CFD2QXL \q0_reg[19]  ( .D(n747), .CP(clk), .CD(n199), .Q(q0[19]) );
  CFD2QXL \q0_reg[20]  ( .D(n748), .CP(clk), .CD(n199), .Q(q0[20]) );
  CFD2QXL \q0_reg[21]  ( .D(n749), .CP(clk), .CD(n199), .Q(q0[21]) );
  CFD2QXL \q0_reg[22]  ( .D(n750), .CP(clk), .CD(n199), .Q(q0[22]) );
  CFD2QXL \q0_reg[23]  ( .D(n751), .CP(clk), .CD(n199), .Q(q0[23]) );
  CFD2QXL \q0_reg[24]  ( .D(n752), .CP(clk), .CD(n199), .Q(q0[24]) );
  CFD2QXL \q0_reg[25]  ( .D(n753), .CP(clk), .CD(n199), .Q(q0[25]) );
  CFD2QXL \q0_reg[26]  ( .D(n754), .CP(clk), .CD(n199), .Q(q0[26]) );
  CFD2QXL \q0_reg[27]  ( .D(n755), .CP(clk), .CD(n199), .Q(q0[27]) );
  CFD2QXL \q0_reg[28]  ( .D(n756), .CP(clk), .CD(n199), .Q(q0[28]) );
  CFD2QXL \q0_reg[29]  ( .D(n757), .CP(clk), .CD(n199), .Q(q0[29]) );
  CFD2QXL \q0_reg[30]  ( .D(n758), .CP(clk), .CD(n199), .Q(q0[30]) );
  CFD2QXL \q0_reg[31]  ( .D(n759), .CP(clk), .CD(n199), .Q(q0[31]) );
  CFD2QXL \cmd0_reg[1]  ( .D(cmd[1]), .CP(clk), .CD(n199), .Q(cmd0[1]) );
  CFD2QXL \cmd0_reg[0]  ( .D(cmd[0]), .CP(clk), .CD(n199), .Q(cmd0[0]) );
  CFD2QXL \cmd1_reg[0]  ( .D(n418), .CP(clk), .CD(n199), .Q(cmd1[0]) );
  CFD2QXL \h0_d_a_reg[1]  ( .D(n605), .CP(clk), .CD(n199), .Q(h0_d_a[1]) );
  CFD2QXL \h0_d_a_reg[2]  ( .D(n606), .CP(clk), .CD(n199), .Q(h0_d_a[2]) );
  CFD2QXL \h0_d_a_reg[4]  ( .D(n607), .CP(clk), .CD(n199), .Q(h0_d_a[4]) );
  CFD2QXL \h0_d_a_reg[5]  ( .D(n608), .CP(clk), .CD(n199), .Q(h0_d_a[5]) );
  CFD2QXL \h0_d_a_reg[6]  ( .D(n609), .CP(clk), .CD(n199), .Q(h0_d_a[6]) );
  CFD2QXL \h0_d_a_reg[0]  ( .D(n610), .CP(clk), .CD(n199), .Q(h0_d_a[0]) );
  CFD2QXL \h0_d_a_reg[3]  ( .D(n611), .CP(clk), .CD(n199), .Q(h0_d_a[3]) );
  CFD2QXL \dout_reg[1]  ( .D(n233), .CP(clk), .CD(n199), .Q(z[1]) );
  CFD2QXL \dout_reg[2]  ( .D(n232), .CP(clk), .CD(n199), .Q(z[2]) );
  CFD2QXL \dout_reg[3]  ( .D(n614), .CP(clk), .CD(n199), .Q(z[3]) );
  CFD2QXL \dout_reg[4]  ( .D(n615), .CP(clk), .CD(n199), .Q(z[4]) );
  CFD2QXL \dout_reg[5]  ( .D(n616), .CP(clk), .CD(n199), .Q(z[5]) );
  CFD2QXL \dout_reg[6]  ( .D(n617), .CP(clk), .CD(n199), .Q(z[6]) );
  CFD2QXL \dout_reg[7]  ( .D(n618), .CP(clk), .CD(n199), .Q(z[7]) );
  CFD2QXL \dout_reg[8]  ( .D(n226), .CP(clk), .CD(n199), .Q(z[8]) );
  CFD2QXL \dout_reg[9]  ( .D(n225), .CP(clk), .CD(n199), .Q(z[9]) );
  CFD2QXL \dout_reg[10]  ( .D(n619), .CP(clk), .CD(n199), .Q(z[10]) );
  CFD2QXL \dout_reg[11]  ( .D(n620), .CP(clk), .CD(n199), .Q(z[11]) );
  CFD2QXL \dout_reg[13]  ( .D(n221), .CP(clk), .CD(n199), .Q(z[13]) );
  CFD2QXL \dout_reg[14]  ( .D(n220), .CP(clk), .CD(n199), .Q(z[14]) );
  CFD2QXL \dout_reg[15]  ( .D(n621), .CP(clk), .CD(n199), .Q(z[15]) );
  CFD2QXL \dout_reg[16]  ( .D(n622), .CP(clk), .CD(n199), .Q(z[16]) );
  CFD2QXL \dout_reg[17]  ( .D(n217), .CP(clk), .CD(n199), .Q(z[17]) );
  CFD2QXL \dout_reg[18]  ( .D(n216), .CP(clk), .CD(n199), .Q(z[18]) );
  CFD2QXL \dout_reg[19]  ( .D(n623), .CP(clk), .CD(n199), .Q(z[19]) );
  CFD2QXL \dout_reg[20]  ( .D(n624), .CP(clk), .CD(n199), .Q(z[20]) );
  CFD2QXL \dout_reg[21]  ( .D(n213), .CP(clk), .CD(n199), .Q(z[21]) );
  CFD2QXL \dout_reg[22]  ( .D(n212), .CP(clk), .CD(n199), .Q(z[22]) );
  CFD2QXL \dout_reg[23]  ( .D(n625), .CP(clk), .CD(n199), .Q(z[23]) );
  CFD2QXL \dout_reg[24]  ( .D(n626), .CP(clk), .CD(n199), .Q(z[24]) );
  CFD2QXL \dout_reg[25]  ( .D(n627), .CP(clk), .CD(n199), .Q(z[25]) );
  CFD2QXL \dout_reg[26]  ( .D(n628), .CP(clk), .CD(n199), .Q(z[26]) );
  CFD2QXL \dout_reg[27]  ( .D(n629), .CP(clk), .CD(n199), .Q(z[27]) );
  CFD2QXL \dout_reg[28]  ( .D(n630), .CP(clk), .CD(n199), .Q(z[28]) );
  CFD2QXL \dout_reg[29]  ( .D(n631), .CP(clk), .CD(n199), .Q(z[29]) );
  CFD2QXL \dout_reg[30]  ( .D(n632), .CP(clk), .CD(n199), .Q(z[30]) );
  CFD2QXL \dout_reg[31]  ( .D(n633), .CP(clk), .CD(n199), .Q(z[31]) );
  CFD2QXL \dout_reg[0]  ( .D(n634), .CP(clk), .CD(n199), .Q(z[0]) );
  CFD2QXL \h0_reg[0]  ( .D(h0_d[0]), .CP(clk), .CD(n199), .Q(h0[0]) );
  CFD2QXL \h0_reg[1]  ( .D(h0_d[1]), .CP(clk), .CD(n199), .Q(h0[1]) );
  CFD2QXL \h0_reg[2]  ( .D(h0_d[2]), .CP(clk), .CD(n199), .Q(h0[2]) );
  CFD2QXL \h0_reg[3]  ( .D(h0_d[3]), .CP(clk), .CD(n199), .Q(h0[3]) );
  CFD2QXL \h0_reg[4]  ( .D(h0_d[4]), .CP(clk), .CD(n199), .Q(h0[4]) );
  CFD2QXL \h0_reg[5]  ( .D(h0_d[5]), .CP(clk), .CD(n199), .Q(h0[5]) );
  CFD2QXL \h0_reg[6]  ( .D(h0_d[6]), .CP(clk), .CD(n199), .Q(h0[6]) );
  CFD2QXL \cmd1_reg[1]  ( .D(n426), .CP(clk), .CD(n199), .Q(cmd1[1]) );
  CFD2QXL \acc_a_reg[63]  ( .D(n298), .CP(clk), .CD(n199), .Q(acc_a[63]) );
  CFD2QXL \acc_a_reg[61]  ( .D(n296), .CP(clk), .CD(n199), .Q(acc_a[61]) );
  CFD2QXL \acc_a_reg[62]  ( .D(n297), .CP(clk), .CD(n199), .Q(acc_a[62]) );
  CFD2QXL \acc_a_reg[60]  ( .D(n295), .CP(clk), .CD(n199), .Q(acc_a[60]) );
  CFD2QXL \acc_a_reg[56]  ( .D(n291), .CP(clk), .CD(n199), .Q(acc_a[56]) );
  CFD2QXL \acc_a_reg[52]  ( .D(n287), .CP(clk), .CD(n199), .Q(acc_a[52]) );
  CMX2XL U297 ( .A0(acc_a[62]), .A1(out[62]), .S(n202), .Z(n297) );
  CMX2XL U287 ( .A0(acc_a[52]), .A1(out[52]), .S(n202), .Z(n287) );
  CMX2XL U291 ( .A0(acc_a[56]), .A1(out[56]), .S(n202), .Z(n291) );
  CMX2XL U298 ( .A0(acc_a[63]), .A1(out[63]), .S(n202), .Z(n298) );
  CMX2XL U295 ( .A0(acc_a[60]), .A1(out[60]), .S(n202), .Z(n295) );
  CMX2XL U296 ( .A0(acc_a[61]), .A1(out[61]), .S(n202), .Z(n296) );
  CND3X1 U234 ( .A(cmd2[0]), .B(cmd2[1]), .C(n1417), .Z(n201) );
  CMX2XL U245 ( .A0(n698), .A1(out[10]), .S(n202), .Z(n245) );
  CMX2XL U288 ( .A0(acc_a[53]), .A1(out[53]), .S(n202), .Z(n288) );
  CMX2XL U235 ( .A0(n690), .A1(out[0]), .S(n202), .Z(n235) );
  CMX2XL U236 ( .A0(n691), .A1(out[1]), .S(n202), .Z(n236) );
  CMX2XL U237 ( .A0(n692), .A1(out[2]), .S(n202), .Z(n237) );
  CMX2XL U238 ( .A0(n693), .A1(out[3]), .S(n202), .Z(n238) );
  CMX2XL U264 ( .A0(acc_a[29]), .A1(out[29]), .S(n202), .Z(n264) );
  CMX2XL U265 ( .A0(acc_a[30]), .A1(out[30]), .S(n202), .Z(n265) );
  CMX2XL U239 ( .A0(n694), .A1(out[4]), .S(n202), .Z(n239) );
  CMX2XL U240 ( .A0(n695), .A1(out[5]), .S(n202), .Z(n240) );
  CMX2XL U241 ( .A0(n696), .A1(out[6]), .S(n202), .Z(n241) );
  CMX2XL U242 ( .A0(n697), .A1(out[7]), .S(n202), .Z(n242) );
  CMX2XL U243 ( .A0(n764), .A1(out[8]), .S(n202), .Z(n243) );
  CMX2XL U244 ( .A0(n762), .A1(out[9]), .S(n202), .Z(n244) );
  CMX2XL U272 ( .A0(acc_a[37]), .A1(out[37]), .S(n202), .Z(n272) );
  CMX2XL U246 ( .A0(n699), .A1(out[11]), .S(n202), .Z(n246) );
  CMX2XL U247 ( .A0(n701), .A1(out[12]), .S(n202), .Z(n247) );
  CMX2XL U248 ( .A0(n767), .A1(out[13]), .S(n202), .Z(n248) );
  CMX2XL U276 ( .A0(acc_a[41]), .A1(out[41]), .S(n202), .Z(n276) );
  CMX2XL U249 ( .A0(n769), .A1(out[14]), .S(n202), .Z(n249) );
  CMX2XL U250 ( .A0(acc_a[15]), .A1(out[15]), .S(n202), .Z(n250) );
  CMX2XL U251 ( .A0(acc_a[16]), .A1(out[16]), .S(n202), .Z(n251) );
  CMX2XL U252 ( .A0(acc_a[17]), .A1(out[17]), .S(n202), .Z(n252) );
  CMX2XL U253 ( .A0(acc_a[18]), .A1(out[18]), .S(n202), .Z(n253) );
  CMX2XL U254 ( .A0(acc_a[19]), .A1(out[19]), .S(n202), .Z(n254) );
  CMX2XL U255 ( .A0(acc_a[20]), .A1(out[20]), .S(n202), .Z(n255) );
  CMX2XL U256 ( .A0(acc_a[21]), .A1(out[21]), .S(n202), .Z(n256) );
  CMX2XL U257 ( .A0(acc_a[22]), .A1(out[22]), .S(n202), .Z(n257) );
  CMX2XL U258 ( .A0(acc_a[23]), .A1(out[23]), .S(n202), .Z(n258) );
  CMX2XL U259 ( .A0(acc_a[24]), .A1(out[24]), .S(n202), .Z(n259) );
  CMX2XL U284 ( .A0(acc_a[49]), .A1(out[49]), .S(n202), .Z(n284) );
  CMX2XL U260 ( .A0(acc_a[25]), .A1(out[25]), .S(n202), .Z(n260) );
  CMX2XL U261 ( .A0(acc_a[26]), .A1(out[26]), .S(n202), .Z(n261) );
  CMX2XL U262 ( .A0(acc_a[27]), .A1(out[27]), .S(n202), .Z(n262) );
  CMX2XL U263 ( .A0(acc_a[28]), .A1(out[28]), .S(n202), .Z(n263) );
  CMX2XL U293 ( .A0(acc_a[58]), .A1(out[58]), .S(n202), .Z(n293) );
  CMX2XL U294 ( .A0(acc_a[59]), .A1(out[59]), .S(n202), .Z(n294) );
  CMX2XL U266 ( .A0(acc_a[31]), .A1(out[31]), .S(n202), .Z(n266) );
  CMX2XL U267 ( .A0(acc_a[32]), .A1(out[32]), .S(n202), .Z(n267) );
  CMX2XL U268 ( .A0(acc_a[33]), .A1(out[33]), .S(n202), .Z(n268) );
  CMX2XL U269 ( .A0(acc_a[34]), .A1(out[34]), .S(n202), .Z(n269) );
  CMX2XL U270 ( .A0(acc_a[35]), .A1(out[35]), .S(n202), .Z(n270) );
  CMX2XL U271 ( .A0(acc_a[36]), .A1(out[36]), .S(n202), .Z(n271) );
  CMX2XL U277 ( .A0(acc_a[42]), .A1(out[42]), .S(n202), .Z(n277) );
  CMX2XL U273 ( .A0(acc_a[38]), .A1(out[38]), .S(n202), .Z(n273) );
  CMX2XL U274 ( .A0(acc_a[39]), .A1(out[39]), .S(n202), .Z(n274) );
  CMX2XL U275 ( .A0(acc_a[40]), .A1(out[40]), .S(n202), .Z(n275) );
  CMX2XL U289 ( .A0(acc_a[54]), .A1(out[54]), .S(n202), .Z(n289) );
  CMX2XL U281 ( .A0(acc_a[46]), .A1(out[46]), .S(n202), .Z(n281) );
  CMX2XL U278 ( .A0(acc_a[43]), .A1(out[43]), .S(n202), .Z(n278) );
  CMX2XL U292 ( .A0(acc_a[57]), .A1(out[57]), .S(n202), .Z(n292) );
  CMX2XL U279 ( .A0(acc_a[44]), .A1(out[44]), .S(n202), .Z(n279) );
  CMX2XL U280 ( .A0(acc_a[45]), .A1(out[45]), .S(n202), .Z(n280) );
  CMX2XL U286 ( .A0(acc_a[51]), .A1(out[51]), .S(n202), .Z(n286) );
  CMX2XL U282 ( .A0(acc_a[47]), .A1(out[47]), .S(n202), .Z(n282) );
  CMX2XL U283 ( .A0(acc_a[48]), .A1(out[48]), .S(n202), .Z(n283) );
  CMX2XL U290 ( .A0(acc_a[55]), .A1(out[55]), .S(n202), .Z(n290) );
  CMX2XL U285 ( .A0(acc_a[50]), .A1(out[50]), .S(n202), .Z(n285) );
  CMX2XL U208 ( .A0(acc[25]), .A1(z[25]), .S(n201), .Z(n209) );
  CMX2XL U207 ( .A0(acc[26]), .A1(z[26]), .S(n201), .Z(n208) );
  CMX2XL U206 ( .A0(acc[27]), .A1(z[27]), .S(n201), .Z(n207) );
  CMX2XL U204 ( .A0(acc[29]), .A1(z[29]), .S(n201), .Z(n205) );
  CMX2XL U205 ( .A0(acc[28]), .A1(z[28]), .S(n201), .Z(n206) );
  CMX2XL U203 ( .A0(acc[30]), .A1(z[30]), .S(n201), .Z(n204) );
  CFD2QX2 \ho_2_reg[1]  ( .D(n636), .CP(clk), .CD(n199), .Q(ho_2[1]) );
  COND1XL \DP_OP_14_298_9081/U360  ( .A(\DP_OP_14_298_9081/n316 ), .B(
        \DP_OP_14_298_9081/n1 ), .C(\DP_OP_14_298_9081/n317 ), .Z(
        \DP_OP_14_298_9081/n315 ) );
  CEOXL \DP_OP_14_298_9081/U316  ( .A(\DP_OP_14_298_9081/n36 ), .B(
        \DP_OP_14_298_9081/n290 ), .Z(\C1/DATA1_32 ) );
  CANR1XL \DP_OP_14_298_9081/U326  ( .A(\DP_OP_14_298_9081/n342 ), .B(
        \DP_OP_14_298_9081/n294 ), .C(\DP_OP_14_298_9081/n295 ), .Z(
        \DP_OP_14_298_9081/n293 ) );
  COND1XL \DP_OP_14_298_9081/U399  ( .A(\DP_OP_14_298_9081/n343 ), .B(
        \DP_OP_14_298_9081/n363 ), .C(\DP_OP_14_298_9081/n344 ), .Z(
        \DP_OP_14_298_9081/n342 ) );
  CANR1X1 \DP_OP_14_298_9081/U463  ( .A(\DP_OP_14_298_9081/n427 ), .B(
        \DP_OP_14_298_9081/n383 ), .C(\DP_OP_14_298_9081/n384 ), .Z(
        \DP_OP_14_298_9081/n1 ) );
  CANR1XL \DP_OP_14_298_9081/U467  ( .A(\DP_OP_14_298_9081/n396 ), .B(
        \DP_OP_14_298_9081/n387 ), .C(\DP_OP_14_298_9081/n388 ), .Z(
        \DP_OP_14_298_9081/n386 ) );
  COND1XL \DP_OP_14_298_9081/U483  ( .A(\DP_OP_14_298_9081/n403 ), .B(
        \DP_OP_14_298_9081/n397 ), .C(\DP_OP_14_298_9081/n398 ), .Z(
        \DP_OP_14_298_9081/n396 ) );
  COND1XL \DP_OP_14_298_9081/U11  ( .A(\DP_OP_14_298_9081/n72 ), .B(
        \DP_OP_14_298_9081/n74 ), .C(\DP_OP_14_298_9081/n73 ), .Z(
        \DP_OP_14_298_9081/n71 ) );
  COND1X1 \DP_OP_14_298_9081/U567  ( .A(\DP_OP_14_298_9081/n455 ), .B(
        \DP_OP_14_298_9081/n451 ), .C(\DP_OP_14_298_9081/n452 ), .Z(
        \DP_OP_14_298_9081/n450 ) );
  CANR1X1 \DP_OP_14_298_9081/U344  ( .A(\DP_OP_14_298_9081/n306 ), .B(
        \DP_OP_14_298_9081/n315 ), .C(\DP_OP_14_298_9081/n307 ), .Z(
        \DP_OP_14_298_9081/n305 ) );
  CEOXL \DP_OP_14_298_9081/U222  ( .A(\DP_OP_14_298_9081/n26 ), .B(
        \DP_OP_14_298_9081/n226 ), .Z(\C1/DATA1_42 ) );
  CEOXL \DP_OP_14_298_9081/U142  ( .A(\DP_OP_14_298_9081/n18 ), .B(
        \DP_OP_14_298_9081/n170 ), .Z(\C1/DATA1_50 ) );
  CANR1X1 \DP_OP_14_298_9081/U295  ( .A(\DP_OP_14_298_9081/n284 ), .B(
        \DP_OP_14_298_9081/n275 ), .C(\DP_OP_14_298_9081/n276 ), .Z(
        \DP_OP_14_298_9081/n270 ) );
  CANR1X1 \DP_OP_14_298_9081/U499  ( .A(\DP_OP_14_298_9081/n420 ), .B(
        \DP_OP_14_298_9081/n407 ), .C(\DP_OP_14_298_9081/n408 ), .Z(
        \DP_OP_14_298_9081/n406 ) );
  CANR1X1 \DP_OP_14_298_9081/U446  ( .A(\DP_OP_14_298_9081/n372 ), .B(
        \DP_OP_14_298_9081/n381 ), .C(\DP_OP_14_298_9081/n373 ), .Z(
        \DP_OP_14_298_9081/n371 ) );
  CANR1X1 \DP_OP_14_298_9081/U171  ( .A(\DP_OP_14_298_9081/n240 ), .B(
        \DP_OP_14_298_9081/n187 ), .C(\DP_OP_14_298_9081/n188 ), .Z(
        \DP_OP_14_298_9081/n3 ) );
  COND1X1 \DP_OP_14_298_9081/U519  ( .A(\DP_OP_14_298_9081/n425 ), .B(
        \DP_OP_14_298_9081/n421 ), .C(\DP_OP_14_298_9081/n422 ), .Z(
        \DP_OP_14_298_9081/n420 ) );
  COND1X1 \DP_OP_14_298_9081/U532  ( .A(\DP_OP_14_298_9081/n428 ), .B(
        \DP_OP_14_298_9081/n448 ), .C(\DP_OP_14_298_9081/n429 ), .Z(
        \DP_OP_14_298_9081/n427 ) );
  CANR1X1 \DP_OP_14_298_9081/U565  ( .A(\DP_OP_14_298_9081/n457 ), .B(
        \DP_OP_14_298_9081/n449 ), .C(\DP_OP_14_298_9081/n450 ), .Z(
        \DP_OP_14_298_9081/n448 ) );
  COND1X1 \DP_OP_14_298_9081/U580  ( .A(\DP_OP_14_298_9081/n461 ), .B(
        \DP_OP_14_298_9081/n458 ), .C(\DP_OP_14_298_9081/n459 ), .Z(
        \DP_OP_14_298_9081/n457 ) );
  CND2X1 \DP_OP_14_298_9081/U559  ( .A(\DP_OP_14_298_9081/n521 ), .B(
        \DP_OP_14_298_9081/n446 ), .Z(\DP_OP_14_298_9081/n64 ) );
  CND2X1 \DP_OP_14_298_9081/U6  ( .A(n1188), .B(\DP_OP_14_298_9081/n70 ), .Z(
        \DP_OP_14_298_9081/n5 ) );
  CND2X1 \DP_OP_14_298_9081/U510  ( .A(\DP_OP_14_298_9081/n515 ), .B(
        \DP_OP_14_298_9081/n415 ), .Z(\DP_OP_14_298_9081/n58 ) );
  CND2X1 \DP_OP_14_298_9081/U484  ( .A(\DP_OP_14_298_9081/n512 ), .B(
        \DP_OP_14_298_9081/n398 ), .Z(\DP_OP_14_298_9081/n55 ) );
  CND2X1 \DP_OP_14_298_9081/U178  ( .A(\DP_OP_14_298_9081/n478 ), .B(
        \DP_OP_14_298_9081/n194 ), .Z(\DP_OP_14_298_9081/n21 ) );
  CND2X1 \DP_OP_14_298_9081/U54  ( .A(\DP_OP_14_298_9081/n466 ), .B(
        \DP_OP_14_298_9081/n106 ), .Z(\DP_OP_14_298_9081/n9 ) );
  CND2X1 \DP_OP_14_298_9081/U236  ( .A(\DP_OP_14_298_9081/n484 ), .B(
        \DP_OP_14_298_9081/n234 ), .Z(\DP_OP_14_298_9081/n27 ) );
  CND2X1 \DP_OP_14_298_9081/U457  ( .A(\DP_OP_14_298_9081/n509 ), .B(
        \DP_OP_14_298_9081/n380 ), .Z(\DP_OP_14_298_9081/n52 ) );
  CND2X1 \DP_OP_14_298_9081/U298  ( .A(\DP_OP_14_298_9081/n490 ), .B(
        \DP_OP_14_298_9081/n278 ), .Z(\DP_OP_14_298_9081/n33 ) );
  CND2X1 \DP_OP_14_298_9081/U218  ( .A(\DP_OP_14_298_9081/n482 ), .B(
        \DP_OP_14_298_9081/n222 ), .Z(\DP_OP_14_298_9081/n25 ) );
  CND2X1 \DP_OP_14_298_9081/U144  ( .A(\DP_OP_14_298_9081/n475 ), .B(
        \DP_OP_14_298_9081/n169 ), .Z(\DP_OP_14_298_9081/n18 ) );
  CNR2X1 \DP_OP_14_298_9081/U44  ( .A(\DP_OP_14_298_9081/n4 ), .B(
        \DP_OP_14_298_9081/n97 ), .Z(\DP_OP_14_298_9081/n95 ) );
  CND2X1 \DP_OP_14_298_9081/U31  ( .A(n1045), .B(acc_a[61]), .Z(
        \DP_OP_14_298_9081/n86 ) );
  CND2X1 \DP_OP_14_298_9081/U57  ( .A(acc[59]), .B(acc_a[59]), .Z(
        \DP_OP_14_298_9081/n106 ) );
  CND2X1 \DP_OP_14_298_9081/U63  ( .A(acc[58]), .B(acc_a[58]), .Z(
        \DP_OP_14_298_9081/n109 ) );
  CND2X1 \DP_OP_14_298_9081/U77  ( .A(n841), .B(acc_a[57]), .Z(
        \DP_OP_14_298_9081/n120 ) );
  CNR2X1 \DP_OP_14_298_9081/U40  ( .A(acc[60]), .B(acc_a[60]), .Z(
        \DP_OP_14_298_9081/n88 ) );
  CND2X1 \DP_OP_14_298_9081/U50  ( .A(\DP_OP_14_298_9081/n115 ), .B(
        \DP_OP_14_298_9081/n103 ), .Z(\DP_OP_14_298_9081/n101 ) );
  CNR2X1 \DP_OP_14_298_9081/U52  ( .A(\DP_OP_14_298_9081/n108 ), .B(
        \DP_OP_14_298_9081/n105 ), .Z(\DP_OP_14_298_9081/n103 ) );
  CNR2X1 \DP_OP_14_298_9081/U56  ( .A(acc[59]), .B(acc_a[59]), .Z(
        \DP_OP_14_298_9081/n105 ) );
  CNR2X1 \DP_OP_14_298_9081/U62  ( .A(acc[58]), .B(acc_a[58]), .Z(
        \DP_OP_14_298_9081/n108 ) );
  CNR2X1 \DP_OP_14_298_9081/U72  ( .A(\DP_OP_14_298_9081/n122 ), .B(
        \DP_OP_14_298_9081/n119 ), .Z(\DP_OP_14_298_9081/n115 ) );
  CNR2X1 \DP_OP_14_298_9081/U76  ( .A(n841), .B(acc_a[57]), .Z(
        \DP_OP_14_298_9081/n119 ) );
  CND2X1 \DP_OP_14_298_9081/U99  ( .A(acc[55]), .B(acc_a[55]), .Z(
        \DP_OP_14_298_9081/n136 ) );
  CND2X1 \DP_OP_14_298_9081/U119  ( .A(acc[53]), .B(acc_a[53]), .Z(
        \DP_OP_14_298_9081/n150 ) );
  CNR2X1 \DP_OP_14_298_9081/U90  ( .A(\DP_OP_14_298_9081/n157 ), .B(
        \DP_OP_14_298_9081/n131 ), .Z(\DP_OP_14_298_9081/n129 ) );
  CND2X1 \DP_OP_14_298_9081/U92  ( .A(\DP_OP_14_298_9081/n145 ), .B(
        \DP_OP_14_298_9081/n133 ), .Z(\DP_OP_14_298_9081/n131 ) );
  CNR2X1 \DP_OP_14_298_9081/U94  ( .A(\DP_OP_14_298_9081/n138 ), .B(
        \DP_OP_14_298_9081/n135 ), .Z(\DP_OP_14_298_9081/n133 ) );
  CNR2X1 \DP_OP_14_298_9081/U98  ( .A(acc[55]), .B(acc_a[55]), .Z(
        \DP_OP_14_298_9081/n135 ) );
  CNR2X1 \DP_OP_14_298_9081/U104  ( .A(acc[54]), .B(acc_a[54]), .Z(
        \DP_OP_14_298_9081/n138 ) );
  CNR2X1 \DP_OP_14_298_9081/U114  ( .A(\DP_OP_14_298_9081/n152 ), .B(
        \DP_OP_14_298_9081/n149 ), .Z(\DP_OP_14_298_9081/n145 ) );
  CNR2X1 \DP_OP_14_298_9081/U118  ( .A(acc[53]), .B(acc_a[53]), .Z(
        \DP_OP_14_298_9081/n149 ) );
  CNR2X1 \DP_OP_14_298_9081/U124  ( .A(acc[52]), .B(acc_a[52]), .Z(
        \DP_OP_14_298_9081/n152 ) );
  CND2X1 \DP_OP_14_298_9081/U134  ( .A(\DP_OP_14_298_9081/n175 ), .B(
        \DP_OP_14_298_9081/n163 ), .Z(\DP_OP_14_298_9081/n157 ) );
  CNR2X1 \DP_OP_14_298_9081/U136  ( .A(\DP_OP_14_298_9081/n168 ), .B(
        \DP_OP_14_298_9081/n165 ), .Z(\DP_OP_14_298_9081/n163 ) );
  CNR2X1 \DP_OP_14_298_9081/U82  ( .A(n1087), .B(acc_a[56]), .Z(
        \DP_OP_14_298_9081/n122 ) );
  CND2X1 \DP_OP_14_298_9081/U138  ( .A(\DP_OP_14_298_9081/n474 ), .B(
        \DP_OP_14_298_9081/n166 ), .Z(\DP_OP_14_298_9081/n17 ) );
  CND2X1 \DP_OP_14_298_9081/U141  ( .A(n1096), .B(acc_a[51]), .Z(
        \DP_OP_14_298_9081/n166 ) );
  CNR2X1 \DP_OP_14_298_9081/U140  ( .A(n1096), .B(acc_a[51]), .Z(
        \DP_OP_14_298_9081/n165 ) );
  CND2X1 \DP_OP_14_298_9081/U147  ( .A(acc[50]), .B(acc_a[50]), .Z(
        \DP_OP_14_298_9081/n169 ) );
  CND2X1 \DP_OP_14_298_9081/U159  ( .A(acc[49]), .B(acc_a[49]), .Z(
        \DP_OP_14_298_9081/n178 ) );
  CND2X1 \DP_OP_14_298_9081/U165  ( .A(acc[48]), .B(acc_a[48]), .Z(
        \DP_OP_14_298_9081/n181 ) );
  CND2X1 \DP_OP_14_298_9081/U181  ( .A(n918), .B(acc_a[47]), .Z(
        \DP_OP_14_298_9081/n194 ) );
  CND2X1 \DP_OP_14_298_9081/U187  ( .A(acc[46]), .B(acc_a[46]), .Z(
        \DP_OP_14_298_9081/n197 ) );
  CND2X1 \DP_OP_14_298_9081/U199  ( .A(n309), .B(acc_a[45]), .Z(
        \DP_OP_14_298_9081/n206 ) );
  CND2X1 \DP_OP_14_298_9081/U205  ( .A(acc[44]), .B(acc_a[44]), .Z(
        \DP_OP_14_298_9081/n209 ) );
  CND2X1 \DP_OP_14_298_9081/U221  ( .A(n917), .B(acc_a[43]), .Z(
        \DP_OP_14_298_9081/n222 ) );
  CND2X1 \DP_OP_14_298_9081/U227  ( .A(acc[42]), .B(acc_a[42]), .Z(
        \DP_OP_14_298_9081/n225 ) );
  CND2X1 \DP_OP_14_298_9081/U239  ( .A(n916), .B(acc_a[41]), .Z(
        \DP_OP_14_298_9081/n234 ) );
  CND2X1 \DP_OP_14_298_9081/U245  ( .A(acc[40]), .B(acc_a[40]), .Z(
        \DP_OP_14_298_9081/n237 ) );
  CND2X1 \DP_OP_14_298_9081/U279  ( .A(n944), .B(acc_a[37]), .Z(
        \DP_OP_14_298_9081/n262 ) );
  CND2X1 \DP_OP_14_298_9081/U285  ( .A(acc[36]), .B(acc_a[36]), .Z(
        \DP_OP_14_298_9081/n265 ) );
  CND2X1 \DP_OP_14_298_9081/U301  ( .A(n915), .B(acc_a[35]), .Z(
        \DP_OP_14_298_9081/n278 ) );
  CND2X1 \DP_OP_14_298_9081/U307  ( .A(acc[34]), .B(acc_a[34]), .Z(
        \DP_OP_14_298_9081/n281 ) );
  CND2X1 \DP_OP_14_298_9081/U315  ( .A(n914), .B(acc_a[33]), .Z(
        \DP_OP_14_298_9081/n286 ) );
  CND2X1 \DP_OP_14_298_9081/U321  ( .A(n913), .B(acc_a[32]), .Z(
        \DP_OP_14_298_9081/n289 ) );
  CND2X1 \DP_OP_14_298_9081/U336  ( .A(acc[31]), .B(acc_a[31]), .Z(
        \DP_OP_14_298_9081/n301 ) );
  CND2X1 \DP_OP_14_298_9081/U342  ( .A(acc[30]), .B(acc_a[30]), .Z(
        \DP_OP_14_298_9081/n304 ) );
  CND2X1 \DP_OP_14_298_9081/U350  ( .A(acc[29]), .B(acc_a[29]), .Z(
        \DP_OP_14_298_9081/n309 ) );
  CND2X1 \DP_OP_14_298_9081/U358  ( .A(acc[28]), .B(acc_a[28]), .Z(
        \DP_OP_14_298_9081/n314 ) );
  CND2X1 \DP_OP_14_298_9081/U372  ( .A(acc[27]), .B(acc_a[27]), .Z(
        \DP_OP_14_298_9081/n325 ) );
  CND2X1 \DP_OP_14_298_9081/U378  ( .A(acc[26]), .B(acc_a[26]), .Z(
        \DP_OP_14_298_9081/n328 ) );
  CND2X1 \DP_OP_14_298_9081/U386  ( .A(acc[25]), .B(acc_a[25]), .Z(
        \DP_OP_14_298_9081/n333 ) );
  CND2X1 \DP_OP_14_298_9081/U392  ( .A(acc[24]), .B(acc_a[24]), .Z(
        \DP_OP_14_298_9081/n336 ) );
  CND2X1 \DP_OP_14_298_9081/U407  ( .A(acc[23]), .B(acc_a[23]), .Z(
        \DP_OP_14_298_9081/n348 ) );
  CND2X1 \DP_OP_14_298_9081/U413  ( .A(n1064), .B(acc_a[22]), .Z(
        \DP_OP_14_298_9081/n351 ) );
  CND2X1 \DP_OP_14_298_9081/U421  ( .A(n1070), .B(acc_a[21]), .Z(
        \DP_OP_14_298_9081/n356 ) );
  CND2X1 \DP_OP_14_298_9081/U427  ( .A(acc[20]), .B(acc_a[20]), .Z(
        \DP_OP_14_298_9081/n359 ) );
  CND2X1 \DP_OP_14_298_9081/U438  ( .A(acc[19]), .B(acc_a[19]), .Z(
        \DP_OP_14_298_9081/n367 ) );
  CND2X1 \DP_OP_14_298_9081/U444  ( .A(n1063), .B(acc_a[18]), .Z(
        \DP_OP_14_298_9081/n370 ) );
  CND2X1 \DP_OP_14_298_9081/U452  ( .A(n1069), .B(acc_a[17]), .Z(
        \DP_OP_14_298_9081/n375 ) );
  CND2X1 \DP_OP_14_298_9081/U460  ( .A(acc[16]), .B(acc_a[16]), .Z(
        \DP_OP_14_298_9081/n380 ) );
  CND2X1 \DP_OP_14_298_9081/U473  ( .A(acc[15]), .B(acc_a[15]), .Z(
        \DP_OP_14_298_9081/n390 ) );
  CND2X1 \DP_OP_14_298_9081/U479  ( .A(n1095), .B(acc_a[14]), .Z(
        \DP_OP_14_298_9081/n393 ) );
  CND2X1 \DP_OP_14_298_9081/U487  ( .A(acc[13]), .B(acc_a[13]), .Z(
        \DP_OP_14_298_9081/n398 ) );
  CND2X1 \DP_OP_14_298_9081/U495  ( .A(acc[12]), .B(acc_a[12]), .Z(
        \DP_OP_14_298_9081/n403 ) );
  CND2X1 \DP_OP_14_298_9081/U505  ( .A(acc[11]), .B(acc_a[11]), .Z(
        \DP_OP_14_298_9081/n410 ) );
  CND2X1 \DP_OP_14_298_9081/U513  ( .A(acc[10]), .B(acc_a[10]), .Z(
        \DP_OP_14_298_9081/n415 ) );
  CND2X1 \DP_OP_14_298_9081/U523  ( .A(acc[9]), .B(acc_a[9]), .Z(
        \DP_OP_14_298_9081/n422 ) );
  CND2X1 \DP_OP_14_298_9081/U529  ( .A(acc[8]), .B(acc_a[8]), .Z(
        \DP_OP_14_298_9081/n425 ) );
  CNR2X1 \DP_OP_14_298_9081/U464  ( .A(\DP_OP_14_298_9081/n405 ), .B(
        \DP_OP_14_298_9081/n385 ), .Z(\DP_OP_14_298_9081/n383 ) );
  CND2X1 \DP_OP_14_298_9081/U466  ( .A(\DP_OP_14_298_9081/n395 ), .B(
        \DP_OP_14_298_9081/n387 ), .Z(\DP_OP_14_298_9081/n385 ) );
  CNR2X1 \DP_OP_14_298_9081/U468  ( .A(\DP_OP_14_298_9081/n392 ), .B(
        \DP_OP_14_298_9081/n389 ), .Z(\DP_OP_14_298_9081/n387 ) );
  CNR2X1 \DP_OP_14_298_9081/U472  ( .A(acc[15]), .B(acc_a[15]), .Z(
        \DP_OP_14_298_9081/n389 ) );
  CNR2X1 \DP_OP_14_298_9081/U482  ( .A(\DP_OP_14_298_9081/n402 ), .B(
        \DP_OP_14_298_9081/n397 ), .Z(\DP_OP_14_298_9081/n395 ) );
  CNR2X1 \DP_OP_14_298_9081/U486  ( .A(acc[13]), .B(acc_a[13]), .Z(
        \DP_OP_14_298_9081/n397 ) );
  CNR2X1 \DP_OP_14_298_9081/U494  ( .A(acc[12]), .B(acc_a[12]), .Z(
        \DP_OP_14_298_9081/n402 ) );
  CND2X1 \DP_OP_14_298_9081/U498  ( .A(\DP_OP_14_298_9081/n419 ), .B(
        \DP_OP_14_298_9081/n407 ), .Z(\DP_OP_14_298_9081/n405 ) );
  CNR2X1 \DP_OP_14_298_9081/U500  ( .A(\DP_OP_14_298_9081/n414 ), .B(
        \DP_OP_14_298_9081/n409 ), .Z(\DP_OP_14_298_9081/n407 ) );
  CNR2X1 \DP_OP_14_298_9081/U504  ( .A(acc[11]), .B(acc_a[11]), .Z(
        \DP_OP_14_298_9081/n409 ) );
  CNR2X1 \DP_OP_14_298_9081/U512  ( .A(acc[10]), .B(acc_a[10]), .Z(
        \DP_OP_14_298_9081/n414 ) );
  CNR2X1 \DP_OP_14_298_9081/U518  ( .A(\DP_OP_14_298_9081/n424 ), .B(
        \DP_OP_14_298_9081/n421 ), .Z(\DP_OP_14_298_9081/n419 ) );
  CNR2X1 \DP_OP_14_298_9081/U522  ( .A(acc[9]), .B(acc_a[9]), .Z(
        \DP_OP_14_298_9081/n421 ) );
  CNR2X1 \DP_OP_14_298_9081/U528  ( .A(acc[8]), .B(acc_a[8]), .Z(
        \DP_OP_14_298_9081/n424 ) );
  CND2X1 \DP_OP_14_298_9081/U540  ( .A(acc[7]), .B(acc_a[7]), .Z(
        \DP_OP_14_298_9081/n433 ) );
  CND2X1 \DP_OP_14_298_9081/U546  ( .A(acc[6]), .B(acc_a[6]), .Z(
        \DP_OP_14_298_9081/n436 ) );
  CND2X1 \DP_OP_14_298_9081/U554  ( .A(acc[5]), .B(acc_a[5]), .Z(
        \DP_OP_14_298_9081/n441 ) );
  CND2X1 \DP_OP_14_298_9081/U562  ( .A(acc[4]), .B(acc_a[4]), .Z(
        \DP_OP_14_298_9081/n446 ) );
  CND2X1 \DP_OP_14_298_9081/U571  ( .A(acc[3]), .B(acc_a[3]), .Z(
        \DP_OP_14_298_9081/n452 ) );
  CND2X1 \DP_OP_14_298_9081/U577  ( .A(acc[2]), .B(acc_a[2]), .Z(
        \DP_OP_14_298_9081/n455 ) );
  CNR2X1 \DP_OP_14_298_9081/U566  ( .A(\DP_OP_14_298_9081/n454 ), .B(
        \DP_OP_14_298_9081/n451 ), .Z(\DP_OP_14_298_9081/n449 ) );
  CNR2X1 \DP_OP_14_298_9081/U570  ( .A(acc[3]), .B(acc_a[3]), .Z(
        \DP_OP_14_298_9081/n451 ) );
  CNR2X1 \DP_OP_14_298_9081/U576  ( .A(acc[2]), .B(acc_a[2]), .Z(
        \DP_OP_14_298_9081/n454 ) );
  CND2X1 \DP_OP_14_298_9081/U584  ( .A(acc[1]), .B(acc_a[1]), .Z(
        \DP_OP_14_298_9081/n459 ) );
  CNR2X1 \DP_OP_14_298_9081/U583  ( .A(acc[1]), .B(acc_a[1]), .Z(
        \DP_OP_14_298_9081/n458 ) );
  CND2X1 \DP_OP_14_298_9081/U589  ( .A(acc[0]), .B(acc_a[0]), .Z(
        \DP_OP_14_298_9081/n461 ) );
  CNR2X1 \DP_OP_14_298_9081/U535  ( .A(\DP_OP_14_298_9081/n435 ), .B(
        \DP_OP_14_298_9081/n432 ), .Z(\DP_OP_14_298_9081/n430 ) );
  CNR2X1 \DP_OP_14_298_9081/U539  ( .A(acc[7]), .B(acc_a[7]), .Z(
        \DP_OP_14_298_9081/n432 ) );
  CNR2X1 \DP_OP_14_298_9081/U545  ( .A(acc[6]), .B(acc_a[6]), .Z(
        \DP_OP_14_298_9081/n435 ) );
  CNR2X1 \DP_OP_14_298_9081/U549  ( .A(\DP_OP_14_298_9081/n445 ), .B(
        \DP_OP_14_298_9081/n440 ), .Z(\DP_OP_14_298_9081/n438 ) );
  CNR2X1 \DP_OP_14_298_9081/U553  ( .A(acc[5]), .B(acc_a[5]), .Z(
        \DP_OP_14_298_9081/n440 ) );
  CNR2X1 \DP_OP_14_298_9081/U561  ( .A(acc[4]), .B(acc_a[4]), .Z(
        \DP_OP_14_298_9081/n445 ) );
  CNR2X1 \DP_OP_14_298_9081/U327  ( .A(\DP_OP_14_298_9081/n320 ), .B(
        \DP_OP_14_298_9081/n296 ), .Z(\DP_OP_14_298_9081/n294 ) );
  CND2X1 \DP_OP_14_298_9081/U329  ( .A(\DP_OP_14_298_9081/n306 ), .B(
        \DP_OP_14_298_9081/n298 ), .Z(\DP_OP_14_298_9081/n296 ) );
  CNR2X1 \DP_OP_14_298_9081/U331  ( .A(\DP_OP_14_298_9081/n303 ), .B(
        \DP_OP_14_298_9081/n300 ), .Z(\DP_OP_14_298_9081/n298 ) );
  CNR2X1 \DP_OP_14_298_9081/U335  ( .A(acc[31]), .B(acc_a[31]), .Z(
        \DP_OP_14_298_9081/n300 ) );
  CNR2X1 \DP_OP_14_298_9081/U341  ( .A(acc[30]), .B(acc_a[30]), .Z(
        \DP_OP_14_298_9081/n303 ) );
  CNR2X1 \DP_OP_14_298_9081/U345  ( .A(\DP_OP_14_298_9081/n313 ), .B(
        \DP_OP_14_298_9081/n308 ), .Z(\DP_OP_14_298_9081/n306 ) );
  CNR2X1 \DP_OP_14_298_9081/U349  ( .A(acc[29]), .B(acc_a[29]), .Z(
        \DP_OP_14_298_9081/n308 ) );
  CNR2X1 \DP_OP_14_298_9081/U357  ( .A(acc[28]), .B(acc_a[28]), .Z(
        \DP_OP_14_298_9081/n313 ) );
  CND2X1 \DP_OP_14_298_9081/U365  ( .A(\DP_OP_14_298_9081/n330 ), .B(
        \DP_OP_14_298_9081/n322 ), .Z(\DP_OP_14_298_9081/n320 ) );
  CNR2X1 \DP_OP_14_298_9081/U367  ( .A(\DP_OP_14_298_9081/n327 ), .B(
        \DP_OP_14_298_9081/n324 ), .Z(\DP_OP_14_298_9081/n322 ) );
  CNR2X1 \DP_OP_14_298_9081/U371  ( .A(acc[27]), .B(acc_a[27]), .Z(
        \DP_OP_14_298_9081/n324 ) );
  CNR2X1 \DP_OP_14_298_9081/U377  ( .A(acc[26]), .B(acc_a[26]), .Z(
        \DP_OP_14_298_9081/n327 ) );
  CNR2X1 \DP_OP_14_298_9081/U381  ( .A(\DP_OP_14_298_9081/n335 ), .B(
        \DP_OP_14_298_9081/n332 ), .Z(\DP_OP_14_298_9081/n330 ) );
  CNR2X1 \DP_OP_14_298_9081/U385  ( .A(acc[25]), .B(acc_a[25]), .Z(
        \DP_OP_14_298_9081/n332 ) );
  CNR2X1 \DP_OP_14_298_9081/U391  ( .A(acc[24]), .B(acc_a[24]), .Z(
        \DP_OP_14_298_9081/n335 ) );
  CNR2X1 \DP_OP_14_298_9081/U398  ( .A(\DP_OP_14_298_9081/n362 ), .B(
        \DP_OP_14_298_9081/n343 ), .Z(\DP_OP_14_298_9081/n341 ) );
  CND2X1 \DP_OP_14_298_9081/U400  ( .A(\DP_OP_14_298_9081/n353 ), .B(
        \DP_OP_14_298_9081/n345 ), .Z(\DP_OP_14_298_9081/n343 ) );
  CNR2X1 \DP_OP_14_298_9081/U402  ( .A(\DP_OP_14_298_9081/n350 ), .B(
        \DP_OP_14_298_9081/n347 ), .Z(\DP_OP_14_298_9081/n345 ) );
  CNR2X1 \DP_OP_14_298_9081/U406  ( .A(acc[23]), .B(acc_a[23]), .Z(
        \DP_OP_14_298_9081/n347 ) );
  CNR2X1 \DP_OP_14_298_9081/U412  ( .A(n1064), .B(acc_a[22]), .Z(
        \DP_OP_14_298_9081/n350 ) );
  CNR2X1 \DP_OP_14_298_9081/U416  ( .A(\DP_OP_14_298_9081/n358 ), .B(
        \DP_OP_14_298_9081/n355 ), .Z(\DP_OP_14_298_9081/n353 ) );
  CNR2X1 \DP_OP_14_298_9081/U420  ( .A(n1070), .B(acc_a[21]), .Z(
        \DP_OP_14_298_9081/n355 ) );
  CNR2X1 \DP_OP_14_298_9081/U426  ( .A(acc[20]), .B(acc_a[20]), .Z(
        \DP_OP_14_298_9081/n358 ) );
  CND2X1 \DP_OP_14_298_9081/U431  ( .A(\DP_OP_14_298_9081/n372 ), .B(
        \DP_OP_14_298_9081/n364 ), .Z(\DP_OP_14_298_9081/n362 ) );
  CNR2X1 \DP_OP_14_298_9081/U433  ( .A(\DP_OP_14_298_9081/n369 ), .B(
        \DP_OP_14_298_9081/n366 ), .Z(\DP_OP_14_298_9081/n364 ) );
  CNR2X1 \DP_OP_14_298_9081/U437  ( .A(acc[19]), .B(acc_a[19]), .Z(
        \DP_OP_14_298_9081/n366 ) );
  CNR2X1 \DP_OP_14_298_9081/U443  ( .A(n1063), .B(acc_a[18]), .Z(
        \DP_OP_14_298_9081/n369 ) );
  CNR2X1 \DP_OP_14_298_9081/U447  ( .A(\DP_OP_14_298_9081/n379 ), .B(
        \DP_OP_14_298_9081/n374 ), .Z(\DP_OP_14_298_9081/n372 ) );
  CNR2X1 \DP_OP_14_298_9081/U451  ( .A(n1069), .B(acc_a[17]), .Z(
        \DP_OP_14_298_9081/n374 ) );
  CNR2X1 \DP_OP_14_298_9081/U459  ( .A(acc[16]), .B(acc_a[16]), .Z(
        \DP_OP_14_298_9081/n379 ) );
  CNR2X1 \DP_OP_14_298_9081/U154  ( .A(\DP_OP_14_298_9081/n180 ), .B(
        \DP_OP_14_298_9081/n177 ), .Z(\DP_OP_14_298_9081/n175 ) );
  CNR2X1 \DP_OP_14_298_9081/U158  ( .A(acc[49]), .B(acc_a[49]), .Z(
        \DP_OP_14_298_9081/n177 ) );
  CNR2X1 \DP_OP_14_298_9081/U164  ( .A(acc[48]), .B(acc_a[48]), .Z(
        \DP_OP_14_298_9081/n180 ) );
  CND2X1 \DP_OP_14_298_9081/U170  ( .A(\DP_OP_14_298_9081/n239 ), .B(
        \DP_OP_14_298_9081/n187 ), .Z(\DP_OP_14_298_9081/n4 ) );
  CNR2X1 \DP_OP_14_298_9081/U172  ( .A(\DP_OP_14_298_9081/n217 ), .B(
        \DP_OP_14_298_9081/n189 ), .Z(\DP_OP_14_298_9081/n187 ) );
  CND2X1 \DP_OP_14_298_9081/U174  ( .A(\DP_OP_14_298_9081/n203 ), .B(
        \DP_OP_14_298_9081/n191 ), .Z(\DP_OP_14_298_9081/n189 ) );
  CNR2X1 \DP_OP_14_298_9081/U176  ( .A(\DP_OP_14_298_9081/n196 ), .B(
        \DP_OP_14_298_9081/n193 ), .Z(\DP_OP_14_298_9081/n191 ) );
  CNR2X1 \DP_OP_14_298_9081/U180  ( .A(n918), .B(acc_a[47]), .Z(
        \DP_OP_14_298_9081/n193 ) );
  CNR2X1 \DP_OP_14_298_9081/U186  ( .A(acc[46]), .B(acc_a[46]), .Z(
        \DP_OP_14_298_9081/n196 ) );
  CNR2X1 \DP_OP_14_298_9081/U194  ( .A(\DP_OP_14_298_9081/n208 ), .B(
        \DP_OP_14_298_9081/n205 ), .Z(\DP_OP_14_298_9081/n203 ) );
  CNR2X1 \DP_OP_14_298_9081/U198  ( .A(n309), .B(acc_a[45]), .Z(
        \DP_OP_14_298_9081/n205 ) );
  CNR2X1 \DP_OP_14_298_9081/U204  ( .A(acc[44]), .B(acc_a[44]), .Z(
        \DP_OP_14_298_9081/n208 ) );
  CND2X1 \DP_OP_14_298_9081/U214  ( .A(\DP_OP_14_298_9081/n231 ), .B(
        \DP_OP_14_298_9081/n219 ), .Z(\DP_OP_14_298_9081/n217 ) );
  CNR2X1 \DP_OP_14_298_9081/U216  ( .A(\DP_OP_14_298_9081/n224 ), .B(
        \DP_OP_14_298_9081/n221 ), .Z(\DP_OP_14_298_9081/n219 ) );
  CNR2X1 \DP_OP_14_298_9081/U220  ( .A(n917), .B(acc_a[43]), .Z(
        \DP_OP_14_298_9081/n221 ) );
  CNR2X1 \DP_OP_14_298_9081/U226  ( .A(acc[42]), .B(acc_a[42]), .Z(
        \DP_OP_14_298_9081/n224 ) );
  CNR2X1 \DP_OP_14_298_9081/U234  ( .A(\DP_OP_14_298_9081/n236 ), .B(
        \DP_OP_14_298_9081/n233 ), .Z(\DP_OP_14_298_9081/n231 ) );
  CNR2X1 \DP_OP_14_298_9081/U238  ( .A(n916), .B(acc_a[41]), .Z(
        \DP_OP_14_298_9081/n233 ) );
  CNR2X1 \DP_OP_14_298_9081/U244  ( .A(acc[40]), .B(acc_a[40]), .Z(
        \DP_OP_14_298_9081/n236 ) );
  CNR2X1 \DP_OP_14_298_9081/U252  ( .A(\DP_OP_14_298_9081/n269 ), .B(
        \DP_OP_14_298_9081/n245 ), .Z(\DP_OP_14_298_9081/n239 ) );
  CND2X1 \DP_OP_14_298_9081/U254  ( .A(\DP_OP_14_298_9081/n259 ), .B(
        \DP_OP_14_298_9081/n247 ), .Z(\DP_OP_14_298_9081/n245 ) );
  CNR2X1 \DP_OP_14_298_9081/U256  ( .A(\DP_OP_14_298_9081/n252 ), .B(
        \DP_OP_14_298_9081/n249 ), .Z(\DP_OP_14_298_9081/n247 ) );
  CNR2X1 \DP_OP_14_298_9081/U260  ( .A(acc[39]), .B(acc_a[39]), .Z(
        \DP_OP_14_298_9081/n249 ) );
  CNR2X1 \DP_OP_14_298_9081/U274  ( .A(\DP_OP_14_298_9081/n264 ), .B(
        \DP_OP_14_298_9081/n261 ), .Z(\DP_OP_14_298_9081/n259 ) );
  CNR2X1 \DP_OP_14_298_9081/U278  ( .A(n944), .B(acc_a[37]), .Z(
        \DP_OP_14_298_9081/n261 ) );
  CNR2X1 \DP_OP_14_298_9081/U284  ( .A(acc[36]), .B(acc_a[36]), .Z(
        \DP_OP_14_298_9081/n264 ) );
  CND2X1 \DP_OP_14_298_9081/U294  ( .A(\DP_OP_14_298_9081/n283 ), .B(
        \DP_OP_14_298_9081/n275 ), .Z(\DP_OP_14_298_9081/n269 ) );
  CNR2X1 \DP_OP_14_298_9081/U296  ( .A(\DP_OP_14_298_9081/n280 ), .B(
        \DP_OP_14_298_9081/n277 ), .Z(\DP_OP_14_298_9081/n275 ) );
  CNR2X1 \DP_OP_14_298_9081/U300  ( .A(n915), .B(acc_a[35]), .Z(
        \DP_OP_14_298_9081/n277 ) );
  CNR2X1 \DP_OP_14_298_9081/U306  ( .A(acc[34]), .B(acc_a[34]), .Z(
        \DP_OP_14_298_9081/n280 ) );
  CNR2X1 \DP_OP_14_298_9081/U310  ( .A(\DP_OP_14_298_9081/n288 ), .B(
        \DP_OP_14_298_9081/n285 ), .Z(\DP_OP_14_298_9081/n283 ) );
  CNR2X1 \DP_OP_14_298_9081/U314  ( .A(n914), .B(acc_a[33]), .Z(
        \DP_OP_14_298_9081/n285 ) );
  CNR2X1 \DP_OP_14_298_9081/U320  ( .A(n913), .B(acc_a[32]), .Z(
        \DP_OP_14_298_9081/n288 ) );
  CNR2X1 \DP_OP_14_298_9081/U146  ( .A(acc[50]), .B(acc_a[50]), .Z(
        \DP_OP_14_298_9081/n168 ) );
  CENX1 \DP_OP_14_298_9081/U563  ( .A(\DP_OP_14_298_9081/n453 ), .B(
        \DP_OP_14_298_9081/n65 ), .Z(\C1/DATA1_3 ) );
  COND1XL \DP_OP_14_298_9081/U573  ( .A(\DP_OP_14_298_9081/n454 ), .B(
        \DP_OP_14_298_9081/n456 ), .C(\DP_OP_14_298_9081/n455 ), .Z(
        \DP_OP_14_298_9081/n453 ) );
  CENX1 \DP_OP_14_298_9081/U555  ( .A(\DP_OP_14_298_9081/n447 ), .B(
        \DP_OP_14_298_9081/n64 ), .Z(\C1/DATA1_4 ) );
  CENX1 \DP_OP_14_298_9081/U5  ( .A(\DP_OP_14_298_9081/n71 ), .B(
        \DP_OP_14_298_9081/n5 ), .Z(\C1/DATA1_63 ) );
  CENX1 \DP_OP_14_298_9081/U506  ( .A(\DP_OP_14_298_9081/n416 ), .B(
        \DP_OP_14_298_9081/n58 ), .Z(\C1/DATA1_10 ) );
  CANR1XL \DP_OP_14_298_9081/U556  ( .A(\DP_OP_14_298_9081/n521 ), .B(
        \DP_OP_14_298_9081/n447 ), .C(\DP_OP_14_298_9081/n444 ), .Z(
        \DP_OP_14_298_9081/n442 ) );
  CENX1 \DP_OP_14_298_9081/U530  ( .A(\DP_OP_14_298_9081/n434 ), .B(
        \DP_OP_14_298_9081/n61 ), .Z(\C1/DATA1_7 ) );
  COND1XL \DP_OP_14_298_9081/U542  ( .A(\DP_OP_14_298_9081/n435 ), .B(
        \DP_OP_14_298_9081/n437 ), .C(\DP_OP_14_298_9081/n436 ), .Z(
        \DP_OP_14_298_9081/n434 ) );
  CANR1XL \DP_OP_14_298_9081/U548  ( .A(\DP_OP_14_298_9081/n438 ), .B(
        \DP_OP_14_298_9081/n447 ), .C(\DP_OP_14_298_9081/n439 ), .Z(
        \DP_OP_14_298_9081/n437 ) );
  CANR1XL \DP_OP_14_298_9081/U380  ( .A(\DP_OP_14_298_9081/n330 ), .B(
        \DP_OP_14_298_9081/n338 ), .C(\DP_OP_14_298_9081/n331 ), .Z(
        \DP_OP_14_298_9081/n329 ) );
  COND1XL \DP_OP_14_298_9081/U395  ( .A(\DP_OP_14_298_9081/n339 ), .B(
        \DP_OP_14_298_9081/n1 ), .C(\DP_OP_14_298_9081/n340 ), .Z(
        \DP_OP_14_298_9081/n338 ) );
  CENX1 \DP_OP_14_298_9081/U166  ( .A(\DP_OP_14_298_9081/n195 ), .B(
        \DP_OP_14_298_9081/n21 ), .Z(\C1/DATA1_47 ) );
  COND1XL \DP_OP_14_298_9081/U183  ( .A(\DP_OP_14_298_9081/n196 ), .B(
        \DP_OP_14_298_9081/n198 ), .C(\DP_OP_14_298_9081/n197 ), .Z(
        \DP_OP_14_298_9081/n195 ) );
  CANR1XL \DP_OP_14_298_9081/U189  ( .A(\DP_OP_14_298_9081/n199 ), .B(
        \DP_OP_14_298_9081/n2 ), .C(\DP_OP_14_298_9081/n200 ), .Z(
        \DP_OP_14_298_9081/n198 ) );
  COND1XL \DP_OP_14_298_9081/U191  ( .A(\DP_OP_14_298_9081/n201 ), .B(
        \DP_OP_14_298_9081/n214 ), .C(\DP_OP_14_298_9081/n202 ), .Z(
        \DP_OP_14_298_9081/n200 ) );
  CANR1XL \DP_OP_14_298_9081/U287  ( .A(\DP_OP_14_298_9081/n267 ), .B(
        \DP_OP_14_298_9081/n2 ), .C(\DP_OP_14_298_9081/n268 ), .Z(
        \DP_OP_14_298_9081/n266 ) );
  COND1XL \DP_OP_14_298_9081/U430  ( .A(\DP_OP_14_298_9081/n362 ), .B(
        \DP_OP_14_298_9081/n1 ), .C(\DP_OP_14_298_9081/n363 ), .Z(
        \DP_OP_14_298_9081/n361 ) );
  CANR1XL \DP_OP_14_298_9081/U352  ( .A(\DP_OP_14_298_9081/n497 ), .B(
        \DP_OP_14_298_9081/n315 ), .C(\DP_OP_14_298_9081/n312 ), .Z(
        \DP_OP_14_298_9081/n310 ) );
  CANR1XL \DP_OP_14_298_9081/U207  ( .A(\DP_OP_14_298_9081/n211 ), .B(
        \DP_OP_14_298_9081/n2 ), .C(\DP_OP_14_298_9081/n212 ), .Z(
        \DP_OP_14_298_9081/n210 ) );
  CANR1XL \DP_OP_14_298_9081/U211  ( .A(\DP_OP_14_298_9081/n215 ), .B(
        \DP_OP_14_298_9081/n240 ), .C(\DP_OP_14_298_9081/n216 ), .Z(
        \DP_OP_14_298_9081/n214 ) );
  CENX1 \DP_OP_14_298_9081/U42  ( .A(\DP_OP_14_298_9081/n107 ), .B(
        \DP_OP_14_298_9081/n9 ), .Z(\C1/DATA1_59 ) );
  COND1XL \DP_OP_14_298_9081/U59  ( .A(\DP_OP_14_298_9081/n108 ), .B(
        \DP_OP_14_298_9081/n110 ), .C(\DP_OP_14_298_9081/n109 ), .Z(
        \DP_OP_14_298_9081/n107 ) );
  CANR1XL \DP_OP_14_298_9081/U65  ( .A(\DP_OP_14_298_9081/n111 ), .B(
        \DP_OP_14_298_9081/n2 ), .C(\DP_OP_14_298_9081/n112 ), .Z(
        \DP_OP_14_298_9081/n110 ) );
  COND1XL \DP_OP_14_298_9081/U67  ( .A(\DP_OP_14_298_9081/n113 ), .B(
        \DP_OP_14_298_9081/n3 ), .C(\DP_OP_14_298_9081/n114 ), .Z(
        \DP_OP_14_298_9081/n112 ) );
  CANR1XL \DP_OP_14_298_9081/U69  ( .A(\DP_OP_14_298_9081/n115 ), .B(
        \DP_OP_14_298_9081/n130 ), .C(\DP_OP_14_298_9081/n118 ), .Z(
        \DP_OP_14_298_9081/n114 ) );
  CENX1 \DP_OP_14_298_9081/U228  ( .A(\DP_OP_14_298_9081/n235 ), .B(
        \DP_OP_14_298_9081/n27 ), .Z(\C1/DATA1_41 ) );
  COND1XL \DP_OP_14_298_9081/U241  ( .A(\DP_OP_14_298_9081/n236 ), .B(
        \DP_OP_14_298_9081/n238 ), .C(\DP_OP_14_298_9081/n237 ), .Z(
        \DP_OP_14_298_9081/n235 ) );
  CANR1XL \DP_OP_14_298_9081/U247  ( .A(\DP_OP_14_298_9081/n239 ), .B(
        \DP_OP_14_298_9081/n2 ), .C(\DP_OP_14_298_9081/n240 ), .Z(
        \DP_OP_14_298_9081/n238 ) );
  CENX1 \DP_OP_14_298_9081/U453  ( .A(\DP_OP_14_298_9081/n381 ), .B(
        \DP_OP_14_298_9081/n52 ), .Z(\C1/DATA1_16 ) );
  CENX1 \DP_OP_14_298_9081/U286  ( .A(\DP_OP_14_298_9081/n279 ), .B(
        \DP_OP_14_298_9081/n33 ), .Z(\C1/DATA1_35 ) );
  COND1XL \DP_OP_14_298_9081/U303  ( .A(\DP_OP_14_298_9081/n280 ), .B(
        \DP_OP_14_298_9081/n282 ), .C(\DP_OP_14_298_9081/n281 ), .Z(
        \DP_OP_14_298_9081/n279 ) );
  CANR1XL \DP_OP_14_298_9081/U309  ( .A(\DP_OP_14_298_9081/n283 ), .B(
        \DP_OP_14_298_9081/n2 ), .C(\DP_OP_14_298_9081/n284 ), .Z(
        \DP_OP_14_298_9081/n282 ) );
  CENX1 \DP_OP_14_298_9081/U206  ( .A(\DP_OP_14_298_9081/n223 ), .B(
        \DP_OP_14_298_9081/n25 ), .Z(\C1/DATA1_43 ) );
  COND1XL \DP_OP_14_298_9081/U223  ( .A(\DP_OP_14_298_9081/n224 ), .B(
        \DP_OP_14_298_9081/n226 ), .C(\DP_OP_14_298_9081/n225 ), .Z(
        \DP_OP_14_298_9081/n223 ) );
  CANR1XL \DP_OP_14_298_9081/U229  ( .A(\DP_OP_14_298_9081/n227 ), .B(
        \DP_OP_14_298_9081/n2 ), .C(\DP_OP_14_298_9081/n228 ), .Z(
        \DP_OP_14_298_9081/n226 ) );
  COND1XL \DP_OP_14_298_9081/U231  ( .A(\DP_OP_14_298_9081/n229 ), .B(
        \DP_OP_14_298_9081/n242 ), .C(\DP_OP_14_298_9081/n230 ), .Z(
        \DP_OP_14_298_9081/n228 ) );
  CANR1XL \DP_OP_14_298_9081/U269  ( .A(\DP_OP_14_298_9081/n255 ), .B(
        \DP_OP_14_298_9081/n2 ), .C(\DP_OP_14_298_9081/n256 ), .Z(
        \DP_OP_14_298_9081/n254 ) );
  COND1XL \DP_OP_14_298_9081/U271  ( .A(\DP_OP_14_298_9081/n257 ), .B(
        \DP_OP_14_298_9081/n270 ), .C(\DP_OP_14_298_9081/n258 ), .Z(
        \DP_OP_14_298_9081/n256 ) );
  CANR1XL \DP_OP_14_298_9081/U127  ( .A(\DP_OP_14_298_9081/n155 ), .B(
        \DP_OP_14_298_9081/n2 ), .C(\DP_OP_14_298_9081/n156 ), .Z(
        \DP_OP_14_298_9081/n154 ) );
  COND1XL \DP_OP_14_298_9081/U129  ( .A(\DP_OP_14_298_9081/n157 ), .B(
        \DP_OP_14_298_9081/n3 ), .C(\DP_OP_14_298_9081/n158 ), .Z(
        \DP_OP_14_298_9081/n156 ) );
  CANR1XL \DP_OP_14_298_9081/U167  ( .A(\DP_OP_14_298_9081/n183 ), .B(
        \DP_OP_14_298_9081/n2 ), .C(\DP_OP_14_298_9081/n184 ), .Z(
        \DP_OP_14_298_9081/n182 ) );
  COND1XL \DP_OP_14_298_9081/U45  ( .A(\DP_OP_14_298_9081/n97 ), .B(
        \DP_OP_14_298_9081/n3 ), .C(\DP_OP_14_298_9081/n98 ), .Z(
        \DP_OP_14_298_9081/n96 ) );
  CANR1XL \DP_OP_14_298_9081/U47  ( .A(\DP_OP_14_298_9081/n99 ), .B(
        \DP_OP_14_298_9081/n130 ), .C(\DP_OP_14_298_9081/n100 ), .Z(
        \DP_OP_14_298_9081/n98 ) );
  CANR1XL \DP_OP_14_298_9081/U362  ( .A(\DP_OP_14_298_9081/n318 ), .B(
        \DP_OP_14_298_9081/n342 ), .C(\DP_OP_14_298_9081/n319 ), .Z(
        \DP_OP_14_298_9081/n317 ) );
  CANR1XL \DP_OP_14_298_9081/U107  ( .A(\DP_OP_14_298_9081/n141 ), .B(
        \DP_OP_14_298_9081/n2 ), .C(\DP_OP_14_298_9081/n142 ), .Z(
        \DP_OP_14_298_9081/n140 ) );
  COND1XL \DP_OP_14_298_9081/U109  ( .A(\DP_OP_14_298_9081/n143 ), .B(
        \DP_OP_14_298_9081/n3 ), .C(\DP_OP_14_298_9081/n144 ), .Z(
        \DP_OP_14_298_9081/n142 ) );
  CANR1XL \DP_OP_14_298_9081/U111  ( .A(\DP_OP_14_298_9081/n145 ), .B(
        \DP_OP_14_298_9081/n160 ), .C(\DP_OP_14_298_9081/n148 ), .Z(
        \DP_OP_14_298_9081/n144 ) );
  CANR1XL \DP_OP_14_298_9081/U17  ( .A(\DP_OP_14_298_9081/n75 ), .B(
        \DP_OP_14_298_9081/n2 ), .C(\DP_OP_14_298_9081/n76 ), .Z(
        \DP_OP_14_298_9081/n74 ) );
  COND1XL \DP_OP_14_298_9081/U19  ( .A(\DP_OP_14_298_9081/n77 ), .B(
        \DP_OP_14_298_9081/n3 ), .C(\DP_OP_14_298_9081/n78 ), .Z(
        \DP_OP_14_298_9081/n76 ) );
  CANR1XL \DP_OP_14_298_9081/U21  ( .A(\DP_OP_14_298_9081/n79 ), .B(
        \DP_OP_14_298_9081/n130 ), .C(\DP_OP_14_298_9081/n80 ), .Z(
        \DP_OP_14_298_9081/n78 ) );
  COND1XL \DP_OP_14_298_9081/U23  ( .A(\DP_OP_14_298_9081/n81 ), .B(
        \DP_OP_14_298_9081/n102 ), .C(\DP_OP_14_298_9081/n82 ), .Z(
        \DP_OP_14_298_9081/n80 ) );
  CANR1XL \DP_OP_14_298_9081/U25  ( .A(\DP_OP_14_298_9081/n91 ), .B(n1190), 
        .C(\DP_OP_14_298_9081/n84 ), .Z(\DP_OP_14_298_9081/n82 ) );
  CANR1XL \DP_OP_14_298_9081/U51  ( .A(\DP_OP_14_298_9081/n118 ), .B(
        \DP_OP_14_298_9081/n103 ), .C(\DP_OP_14_298_9081/n104 ), .Z(
        \DP_OP_14_298_9081/n102 ) );
  COND1XL \DP_OP_14_298_9081/U53  ( .A(\DP_OP_14_298_9081/n109 ), .B(
        \DP_OP_14_298_9081/n105 ), .C(\DP_OP_14_298_9081/n106 ), .Z(
        \DP_OP_14_298_9081/n104 ) );
  COND1XL \DP_OP_14_298_9081/U73  ( .A(\DP_OP_14_298_9081/n123 ), .B(
        \DP_OP_14_298_9081/n119 ), .C(\DP_OP_14_298_9081/n120 ), .Z(
        \DP_OP_14_298_9081/n118 ) );
  CANR1XL \DP_OP_14_298_9081/U85  ( .A(\DP_OP_14_298_9081/n125 ), .B(
        \DP_OP_14_298_9081/n2 ), .C(\DP_OP_14_298_9081/n126 ), .Z(
        \DP_OP_14_298_9081/n124 ) );
  COND1XL \DP_OP_14_298_9081/U87  ( .A(\DP_OP_14_298_9081/n127 ), .B(
        \DP_OP_14_298_9081/n3 ), .C(\DP_OP_14_298_9081/n128 ), .Z(
        \DP_OP_14_298_9081/n126 ) );
  CANR1XL \DP_OP_14_298_9081/U93  ( .A(\DP_OP_14_298_9081/n148 ), .B(
        \DP_OP_14_298_9081/n133 ), .C(\DP_OP_14_298_9081/n134 ), .Z(
        \DP_OP_14_298_9081/n132 ) );
  COND1XL \DP_OP_14_298_9081/U95  ( .A(\DP_OP_14_298_9081/n139 ), .B(
        \DP_OP_14_298_9081/n135 ), .C(\DP_OP_14_298_9081/n136 ), .Z(
        \DP_OP_14_298_9081/n134 ) );
  COND1XL \DP_OP_14_298_9081/U115  ( .A(\DP_OP_14_298_9081/n153 ), .B(
        \DP_OP_14_298_9081/n149 ), .C(\DP_OP_14_298_9081/n150 ), .Z(
        \DP_OP_14_298_9081/n148 ) );
  COND1XL \DP_OP_14_298_9081/U137  ( .A(\DP_OP_14_298_9081/n169 ), .B(
        \DP_OP_14_298_9081/n165 ), .C(\DP_OP_14_298_9081/n166 ), .Z(
        \DP_OP_14_298_9081/n164 ) );
  CENX1 \DP_OP_14_298_9081/U126  ( .A(\DP_OP_14_298_9081/n167 ), .B(
        \DP_OP_14_298_9081/n17 ), .Z(\C1/DATA1_51 ) );
  COND1XL \DP_OP_14_298_9081/U143  ( .A(\DP_OP_14_298_9081/n168 ), .B(
        \DP_OP_14_298_9081/n170 ), .C(\DP_OP_14_298_9081/n169 ), .Z(
        \DP_OP_14_298_9081/n167 ) );
  CANR1XL \DP_OP_14_298_9081/U149  ( .A(\DP_OP_14_298_9081/n171 ), .B(
        \DP_OP_14_298_9081/n2 ), .C(\DP_OP_14_298_9081/n172 ), .Z(
        \DP_OP_14_298_9081/n170 ) );
  COND1XL \DP_OP_14_298_9081/U151  ( .A(\DP_OP_14_298_9081/n173 ), .B(
        \DP_OP_14_298_9081/n3 ), .C(\DP_OP_14_298_9081/n174 ), .Z(
        \DP_OP_14_298_9081/n172 ) );
  COND1XL \DP_OP_14_298_9081/U155  ( .A(\DP_OP_14_298_9081/n181 ), .B(
        \DP_OP_14_298_9081/n177 ), .C(\DP_OP_14_298_9081/n178 ), .Z(
        \DP_OP_14_298_9081/n176 ) );
  COND1XL \DP_OP_14_298_9081/U173  ( .A(\DP_OP_14_298_9081/n189 ), .B(
        \DP_OP_14_298_9081/n218 ), .C(\DP_OP_14_298_9081/n190 ), .Z(
        \DP_OP_14_298_9081/n188 ) );
  CANR1XL \DP_OP_14_298_9081/U175  ( .A(\DP_OP_14_298_9081/n204 ), .B(
        \DP_OP_14_298_9081/n191 ), .C(\DP_OP_14_298_9081/n192 ), .Z(
        \DP_OP_14_298_9081/n190 ) );
  COND1XL \DP_OP_14_298_9081/U177  ( .A(\DP_OP_14_298_9081/n197 ), .B(
        \DP_OP_14_298_9081/n193 ), .C(\DP_OP_14_298_9081/n194 ), .Z(
        \DP_OP_14_298_9081/n192 ) );
  COND1XL \DP_OP_14_298_9081/U195  ( .A(\DP_OP_14_298_9081/n209 ), .B(
        \DP_OP_14_298_9081/n205 ), .C(\DP_OP_14_298_9081/n206 ), .Z(
        \DP_OP_14_298_9081/n204 ) );
  CANR1XL \DP_OP_14_298_9081/U215  ( .A(\DP_OP_14_298_9081/n232 ), .B(
        \DP_OP_14_298_9081/n219 ), .C(\DP_OP_14_298_9081/n220 ), .Z(
        \DP_OP_14_298_9081/n218 ) );
  COND1XL \DP_OP_14_298_9081/U217  ( .A(\DP_OP_14_298_9081/n225 ), .B(
        \DP_OP_14_298_9081/n221 ), .C(\DP_OP_14_298_9081/n222 ), .Z(
        \DP_OP_14_298_9081/n220 ) );
  COND1XL \DP_OP_14_298_9081/U235  ( .A(\DP_OP_14_298_9081/n237 ), .B(
        \DP_OP_14_298_9081/n233 ), .C(\DP_OP_14_298_9081/n234 ), .Z(
        \DP_OP_14_298_9081/n232 ) );
  CANR1XL \DP_OP_14_298_9081/U255  ( .A(\DP_OP_14_298_9081/n260 ), .B(
        \DP_OP_14_298_9081/n247 ), .C(\DP_OP_14_298_9081/n248 ), .Z(
        \DP_OP_14_298_9081/n246 ) );
  COND1XL \DP_OP_14_298_9081/U257  ( .A(\DP_OP_14_298_9081/n253 ), .B(
        \DP_OP_14_298_9081/n249 ), .C(\DP_OP_14_298_9081/n250 ), .Z(
        \DP_OP_14_298_9081/n248 ) );
  COND1XL \DP_OP_14_298_9081/U275  ( .A(\DP_OP_14_298_9081/n265 ), .B(
        \DP_OP_14_298_9081/n261 ), .C(\DP_OP_14_298_9081/n262 ), .Z(
        \DP_OP_14_298_9081/n260 ) );
  COND1XL \DP_OP_14_298_9081/U297  ( .A(\DP_OP_14_298_9081/n281 ), .B(
        \DP_OP_14_298_9081/n277 ), .C(\DP_OP_14_298_9081/n278 ), .Z(
        \DP_OP_14_298_9081/n276 ) );
  COND1XL \DP_OP_14_298_9081/U311  ( .A(\DP_OP_14_298_9081/n289 ), .B(
        \DP_OP_14_298_9081/n285 ), .C(\DP_OP_14_298_9081/n286 ), .Z(
        \DP_OP_14_298_9081/n284 ) );
  COND1XL \DP_OP_14_298_9081/U328  ( .A(\DP_OP_14_298_9081/n296 ), .B(
        \DP_OP_14_298_9081/n321 ), .C(\DP_OP_14_298_9081/n297 ), .Z(
        \DP_OP_14_298_9081/n295 ) );
  CANR1XL \DP_OP_14_298_9081/U330  ( .A(\DP_OP_14_298_9081/n307 ), .B(
        \DP_OP_14_298_9081/n298 ), .C(\DP_OP_14_298_9081/n299 ), .Z(
        \DP_OP_14_298_9081/n297 ) );
  COND1XL \DP_OP_14_298_9081/U332  ( .A(\DP_OP_14_298_9081/n304 ), .B(
        \DP_OP_14_298_9081/n300 ), .C(\DP_OP_14_298_9081/n301 ), .Z(
        \DP_OP_14_298_9081/n299 ) );
  COND1XL \DP_OP_14_298_9081/U346  ( .A(\DP_OP_14_298_9081/n314 ), .B(
        \DP_OP_14_298_9081/n308 ), .C(\DP_OP_14_298_9081/n309 ), .Z(
        \DP_OP_14_298_9081/n307 ) );
  CANR1XL \DP_OP_14_298_9081/U366  ( .A(\DP_OP_14_298_9081/n331 ), .B(
        \DP_OP_14_298_9081/n322 ), .C(\DP_OP_14_298_9081/n323 ), .Z(
        \DP_OP_14_298_9081/n321 ) );
  COND1XL \DP_OP_14_298_9081/U368  ( .A(\DP_OP_14_298_9081/n328 ), .B(
        \DP_OP_14_298_9081/n324 ), .C(\DP_OP_14_298_9081/n325 ), .Z(
        \DP_OP_14_298_9081/n323 ) );
  COND1XL \DP_OP_14_298_9081/U382  ( .A(\DP_OP_14_298_9081/n336 ), .B(
        \DP_OP_14_298_9081/n332 ), .C(\DP_OP_14_298_9081/n333 ), .Z(
        \DP_OP_14_298_9081/n331 ) );
  CANR1XL \DP_OP_14_298_9081/U401  ( .A(\DP_OP_14_298_9081/n354 ), .B(
        \DP_OP_14_298_9081/n345 ), .C(\DP_OP_14_298_9081/n346 ), .Z(
        \DP_OP_14_298_9081/n344 ) );
  COND1XL \DP_OP_14_298_9081/U403  ( .A(\DP_OP_14_298_9081/n351 ), .B(
        \DP_OP_14_298_9081/n347 ), .C(\DP_OP_14_298_9081/n348 ), .Z(
        \DP_OP_14_298_9081/n346 ) );
  COND1XL \DP_OP_14_298_9081/U417  ( .A(\DP_OP_14_298_9081/n359 ), .B(
        \DP_OP_14_298_9081/n355 ), .C(\DP_OP_14_298_9081/n356 ), .Z(
        \DP_OP_14_298_9081/n354 ) );
  CANR1XL \DP_OP_14_298_9081/U432  ( .A(\DP_OP_14_298_9081/n373 ), .B(
        \DP_OP_14_298_9081/n364 ), .C(\DP_OP_14_298_9081/n365 ), .Z(
        \DP_OP_14_298_9081/n363 ) );
  COND1XL \DP_OP_14_298_9081/U434  ( .A(\DP_OP_14_298_9081/n370 ), .B(
        \DP_OP_14_298_9081/n366 ), .C(\DP_OP_14_298_9081/n367 ), .Z(
        \DP_OP_14_298_9081/n365 ) );
  COND1XL \DP_OP_14_298_9081/U448  ( .A(\DP_OP_14_298_9081/n380 ), .B(
        \DP_OP_14_298_9081/n374 ), .C(\DP_OP_14_298_9081/n375 ), .Z(
        \DP_OP_14_298_9081/n373 ) );
  COND1XL \DP_OP_14_298_9081/U469  ( .A(\DP_OP_14_298_9081/n393 ), .B(
        \DP_OP_14_298_9081/n389 ), .C(\DP_OP_14_298_9081/n390 ), .Z(
        \DP_OP_14_298_9081/n388 ) );
  COND1XL \DP_OP_14_298_9081/U501  ( .A(\DP_OP_14_298_9081/n415 ), .B(
        \DP_OP_14_298_9081/n409 ), .C(\DP_OP_14_298_9081/n410 ), .Z(
        \DP_OP_14_298_9081/n408 ) );
  CANR1XL \DP_OP_14_298_9081/U534  ( .A(\DP_OP_14_298_9081/n439 ), .B(
        \DP_OP_14_298_9081/n430 ), .C(\DP_OP_14_298_9081/n431 ), .Z(
        \DP_OP_14_298_9081/n429 ) );
  COND1XL \DP_OP_14_298_9081/U536  ( .A(\DP_OP_14_298_9081/n436 ), .B(
        \DP_OP_14_298_9081/n432 ), .C(\DP_OP_14_298_9081/n433 ), .Z(
        \DP_OP_14_298_9081/n431 ) );
  COND1XL \DP_OP_14_298_9081/U550  ( .A(\DP_OP_14_298_9081/n446 ), .B(
        \DP_OP_14_298_9081/n440 ), .C(\DP_OP_14_298_9081/n441 ), .Z(
        \DP_OP_14_298_9081/n439 ) );
  CFD2QX2 \acc_reg[24]  ( .D(n172), .CP(clk), .CD(n199), .Q(acc[24]) );
  CFD2QX2 \acc_reg[23]  ( .D(n173), .CP(clk), .CD(n199), .Q(acc[23]) );
  CFD2QX2 \acc_reg[15]  ( .D(n181), .CP(clk), .CD(n199), .Q(acc[15]) );
  CFD2QX2 \acc_reg[16]  ( .D(n180), .CP(clk), .CD(n199), .Q(acc[16]) );
  CFD2QX2 \acc_reg[9]  ( .D(n187), .CP(clk), .CD(n199), .Q(acc[9]) );
  CFD2QX2 \acc_reg[8]  ( .D(n188), .CP(clk), .CD(n199), .Q(acc[8]) );
  CFD2QX2 \acc_reg[13]  ( .D(n183), .CP(clk), .CD(n199), .Q(acc[13]) );
  CFD2QX2 \acc_reg[36]  ( .D(n160), .CP(clk), .CD(n199), .Q(acc[36]) );
  CEOXL \DP_OP_14_298_9081/U262  ( .A(\DP_OP_14_298_9081/n30 ), .B(
        \DP_OP_14_298_9081/n254 ), .Z(\C1/DATA1_38 ) );
  CENX1 \DP_OP_14_298_9081/U64  ( .A(\DP_OP_14_298_9081/n121 ), .B(
        \DP_OP_14_298_9081/n11 ), .Z(\C1/DATA1_57 ) );
  COND1XL \DP_OP_14_298_9081/U79  ( .A(\DP_OP_14_298_9081/n122 ), .B(
        \DP_OP_14_298_9081/n124 ), .C(\DP_OP_14_298_9081/n123 ), .Z(
        \DP_OP_14_298_9081/n121 ) );
  CND2X1 \DP_OP_14_298_9081/U74  ( .A(\DP_OP_14_298_9081/n468 ), .B(
        \DP_OP_14_298_9081/n120 ), .Z(\DP_OP_14_298_9081/n11 ) );
  CEOXL \DP_OP_14_298_9081/U120  ( .A(\DP_OP_14_298_9081/n16 ), .B(
        \DP_OP_14_298_9081/n154 ), .Z(\C1/DATA1_52 ) );
  CFD2X2 \acc_reg[51]  ( .D(n145), .CP(clk), .CD(n199), .Q(n1096) );
  CFD2X1 \acc_reg[56]  ( .D(n140), .CP(clk), .CD(n199), .Q(n1087) );
  CFD2X1 \acc_reg[21]  ( .D(n175), .CP(clk), .CD(n199), .Q(n1070) );
  CFD2X1 \acc_reg[17]  ( .D(n179), .CP(clk), .CD(n199), .Q(n1069) );
  CFD2X1 \acc_reg[22]  ( .D(n174), .CP(clk), .CD(n199), .Q(n1064) );
  CFD2X1 \acc_reg[18]  ( .D(n178), .CP(clk), .CD(n199), .Q(n1063) );
  CENX1 \DP_OP_14_298_9081/U84  ( .A(\DP_OP_14_298_9081/n137 ), .B(
        \DP_OP_14_298_9081/n13 ), .Z(\C1/DATA1_55 ) );
  COND1XL \DP_OP_14_298_9081/U101  ( .A(\DP_OP_14_298_9081/n138 ), .B(
        \DP_OP_14_298_9081/n140 ), .C(\DP_OP_14_298_9081/n139 ), .Z(
        \DP_OP_14_298_9081/n137 ) );
  CND2X1 \DP_OP_14_298_9081/U96  ( .A(\DP_OP_14_298_9081/n470 ), .B(
        \DP_OP_14_298_9081/n136 ), .Z(\DP_OP_14_298_9081/n13 ) );
  CEOXL \DP_OP_14_298_9081/U10  ( .A(\DP_OP_14_298_9081/n6 ), .B(
        \DP_OP_14_298_9081/n74 ), .Z(\C1/DATA1_62 ) );
  CEOXL \DP_OP_14_298_9081/U240  ( .A(\DP_OP_14_298_9081/n28 ), .B(
        \DP_OP_14_298_9081/n238 ), .Z(\C1/DATA1_40 ) );
  CFD2X1 \acc_reg[61]  ( .D(n135), .CP(clk), .CD(n199), .Q(n1045) );
  CFD2X1 \acc_reg[37]  ( .D(n159), .CP(clk), .CD(n199), .Q(n944) );
  CFD4X2 \ho_2_reg[0]  ( .D(n931), .CP(clk), .SD(n199), .Q(n921), .QN(ho_2[0])
         );
  CFD2X2 \acc_reg[55]  ( .D(n141), .CP(clk), .CD(n199), .Q(acc[55]) );
  CFD2QX2 \ho_2_reg[2]  ( .D(n637), .CP(clk), .CD(n199), .Q(ho_2[2]) );
  CFD2XL \acc_reg[62]  ( .D(n134), .CP(clk), .CD(n199), .Q(n925), .QN(n924) );
  CFD2QX2 \acc_reg[40]  ( .D(n156), .CP(clk), .CD(n199), .Q(acc[40]) );
  CFD2X1 \acc_reg[47]  ( .D(n149), .CP(clk), .CD(n199), .Q(n918) );
  CFD2X1 \acc_reg[43]  ( .D(n153), .CP(clk), .CD(n199), .Q(n917) );
  CFD2X1 \acc_reg[41]  ( .D(n155), .CP(clk), .CD(n199), .Q(n916) );
  CFD2X1 \acc_reg[35]  ( .D(n161), .CP(clk), .CD(n199), .Q(n915) );
  CFD2X1 \acc_reg[33]  ( .D(n163), .CP(clk), .CD(n199), .Q(n914) );
  CFD2X1 \acc_reg[32]  ( .D(n164), .CP(clk), .CD(n199), .Q(n913) );
  CEOXL \DP_OP_14_298_9081/U200  ( .A(\DP_OP_14_298_9081/n24 ), .B(
        \DP_OP_14_298_9081/n210 ), .Z(\C1/DATA1_44 ) );
  CFD2X2 \acc_reg[44]  ( .D(n152), .CP(clk), .CD(n199), .Q(acc[44]) );
  CFD2X2 \acc_reg[49]  ( .D(n147), .CP(clk), .CD(n199), .Q(acc[49]) );
  CFD2QX2 \acc_reg[59]  ( .D(n137), .CP(clk), .CD(n199), .Q(acc[59]) );
  CEOXL \DP_OP_14_298_9081/U58  ( .A(\DP_OP_14_298_9081/n10 ), .B(
        \DP_OP_14_298_9081/n110 ), .Z(\C1/DATA1_58 ) );
  CND2X1 \DP_OP_14_298_9081/U60  ( .A(\DP_OP_14_298_9081/n467 ), .B(
        \DP_OP_14_298_9081/n109 ), .Z(\DP_OP_14_298_9081/n10 ) );
  CFD2X1 \acc_reg[58]  ( .D(n138), .CP(clk), .CD(n199), .Q(acc[58]) );
  CFD2X2 \acc_reg[53]  ( .D(n143), .CP(clk), .CD(n199), .Q(acc[53]) );
  CFD2X2 \acc_reg[60]  ( .D(n136), .CP(clk), .CD(n199), .Q(acc[60]) );
  CFD2X1 \acc_reg[57]  ( .D(n139), .CP(clk), .CD(n199), .Q(n841) );
  CFD2QX4 \acc_reg[50]  ( .D(n146), .CP(clk), .CD(n199), .Q(acc[50]) );
  COND1XL \DP_OP_14_298_9081/U121  ( .A(\DP_OP_14_298_9081/n152 ), .B(
        \DP_OP_14_298_9081/n154 ), .C(\DP_OP_14_298_9081/n153 ), .Z(
        \DP_OP_14_298_9081/n151 ) );
  CND2X1 \DP_OP_14_298_9081/U116  ( .A(\DP_OP_14_298_9081/n472 ), .B(
        \DP_OP_14_298_9081/n150 ), .Z(\DP_OP_14_298_9081/n15 ) );
  CEOXL \DP_OP_14_298_9081/U32  ( .A(\DP_OP_14_298_9081/n8 ), .B(
        \DP_OP_14_298_9081/n94 ), .Z(\C1/DATA1_60 ) );
  CFD2QX2 \acc_reg[52]  ( .D(n144), .CP(clk), .CD(n199), .Q(acc[52]) );
  CFD2QX2 \acc_reg[19]  ( .D(n177), .CP(clk), .CD(n199), .Q(acc[19]) );
  CEOXL \DP_OP_14_298_9081/U160  ( .A(\DP_OP_14_298_9081/n20 ), .B(
        \DP_OP_14_298_9081/n182 ), .Z(\C1/DATA1_48 ) );
  CENX1 \DP_OP_14_298_9081/U148  ( .A(\DP_OP_14_298_9081/n179 ), .B(
        \DP_OP_14_298_9081/n19 ), .Z(\C1/DATA1_49 ) );
  COND1XL \DP_OP_14_298_9081/U161  ( .A(\DP_OP_14_298_9081/n180 ), .B(
        \DP_OP_14_298_9081/n182 ), .C(\DP_OP_14_298_9081/n181 ), .Z(
        \DP_OP_14_298_9081/n179 ) );
  CND2X1 \DP_OP_14_298_9081/U156  ( .A(\DP_OP_14_298_9081/n476 ), .B(
        \DP_OP_14_298_9081/n178 ), .Z(\DP_OP_14_298_9081/n19 ) );
  CAOR2XL U304 ( .A(pushin), .B(h[28]), .C(n1432), .D(h0[28]), .Z(h0_d[28]) );
  CAOR2XL U306 ( .A(pushin), .B(h[26]), .C(n1431), .D(h0[26]), .Z(h0_d[26]) );
  CAOR2XL U316 ( .A(pushin), .B(h[16]), .C(n1430), .D(h0[16]), .Z(h0_d[16]) );
  CAOR2XL U303 ( .A(pushin), .B(h[29]), .C(n1431), .D(h0[29]), .Z(h0_d[29]) );
  CAOR2XL U317 ( .A(pushin), .B(h[15]), .C(n1431), .D(h0[15]), .Z(h0_d[15]) );
  CAOR2XL U307 ( .A(pushin), .B(h[25]), .C(n1432), .D(h0[25]), .Z(h0_d[25]) );
  CAOR2XL U315 ( .A(pushin), .B(h[17]), .C(n1431), .D(h0[17]), .Z(h0_d[17]) );
  CAOR2XL U301 ( .A(pushin), .B(h[31]), .C(n1430), .D(h0[31]), .Z(h0_d[31]) );
  CAOR2XL U314 ( .A(pushin), .B(h[18]), .C(n1432), .D(h0[18]), .Z(h0_d[18]) );
  CAOR2XL U308 ( .A(pushin), .B(h[24]), .C(n1430), .D(h0[24]), .Z(h0_d[24]) );
  CAOR2XL U313 ( .A(pushin), .B(h[19]), .C(n1432), .D(h0[19]), .Z(h0_d[19]) );
  CAOR2XL U312 ( .A(pushin), .B(h[20]), .C(n1432), .D(h0[20]), .Z(h0_d[20]) );
  CAOR2XL U311 ( .A(pushin), .B(h[21]), .C(n1430), .D(h0[21]), .Z(h0_d[21]) );
  CAOR2XL U360 ( .A(pushin), .B(q[4]), .C(n1432), .D(q0[4]), .Z(q0_d[4]) );
  CAOR2XL U309 ( .A(pushin), .B(h[23]), .C(n1431), .D(h0[23]), .Z(h0_d[23]) );
  CAOR2XL U359 ( .A(pushin), .B(q[5]), .C(n1431), .D(q0[5]), .Z(q0_d[5]) );
  CAOR2XL U310 ( .A(pushin), .B(h[22]), .C(n1430), .D(h0[22]), .Z(h0_d[22]) );
  CAOR2XL U356 ( .A(pushin), .B(q[8]), .C(n1431), .D(q0[8]), .Z(q0_d[8]) );
  CAOR2XL U358 ( .A(pushin), .B(q[6]), .C(n1432), .D(q0[6]), .Z(q0_d[6]) );
  CAOR2XL U357 ( .A(pushin), .B(q[7]), .C(n1430), .D(q0[7]), .Z(q0_d[7]) );
  CAOR2XL U323 ( .A(pushin), .B(h[9]), .C(n1431), .D(h0[9]), .Z(h0_d[9]) );
  CND2XL \DP_OP_14_298_9081/U9  ( .A(acc[63]), .B(acc_a[63]), .Z(
        \DP_OP_14_298_9081/n70 ) );
  CAOR2XL U324 ( .A(pushin), .B(h[8]), .C(n1431), .D(h0[8]), .Z(h0_d[8]) );
  CAOR2XL U318 ( .A(pushin), .B(h[14]), .C(n1432), .D(h0[14]), .Z(h0_d[14]) );
  CAOR2XL U340 ( .A(pushin), .B(q[24]), .C(n1430), .D(q0[24]), .Z(q0_d[24]) );
  CAOR2XL U338 ( .A(pushin), .B(q[26]), .C(n1432), .D(q0[26]), .Z(q0_d[26]) );
  CAOR2XL U337 ( .A(pushin), .B(q[27]), .C(n1432), .D(q0[27]), .Z(q0_d[27]) );
  CAOR2XL U322 ( .A(pushin), .B(h[10]), .C(n1431), .D(h0[10]), .Z(h0_d[10]) );
  CAOR2XL U321 ( .A(pushin), .B(h[11]), .C(n1430), .D(h0[11]), .Z(h0_d[11]) );
  CAOR2XL U325 ( .A(pushin), .B(h[7]), .C(n1430), .D(h0[7]), .Z(h0_d[7]) );
  CAOR2XL U339 ( .A(pushin), .B(q[25]), .C(n1431), .D(q0[25]), .Z(q0_d[25]) );
  CAOR2XL U336 ( .A(pushin), .B(q[28]), .C(n1431), .D(q0[28]), .Z(q0_d[28]) );
  CAOR2XL U335 ( .A(pushin), .B(q[29]), .C(n1430), .D(q0[29]), .Z(q0_d[29]) );
  CAOR2XL U334 ( .A(pushin), .B(q[30]), .C(n1430), .D(q0[30]), .Z(q0_d[30]) );
  CAOR2XL U333 ( .A(pushin), .B(q[31]), .C(n1430), .D(q0[31]), .Z(q0_d[31]) );
  CAOR2XL U364 ( .A(pushin), .B(q[0]), .C(n1432), .D(q0[0]), .Z(q0_d[0]) );
  CAOR2XL U348 ( .A(pushin), .B(q[16]), .C(n1430), .D(q0[16]), .Z(q0_d[16]) );
  CAOR2XL U347 ( .A(pushin), .B(q[17]), .C(n1430), .D(q0[17]), .Z(q0_d[17]) );
  CAOR2XL U346 ( .A(pushin), .B(q[18]), .C(n1432), .D(q0[18]), .Z(q0_d[18]) );
  CAOR2XL U345 ( .A(pushin), .B(q[19]), .C(n1432), .D(q0[19]), .Z(q0_d[19]) );
  CAOR2XL U344 ( .A(pushin), .B(q[20]), .C(n1430), .D(q0[20]), .Z(q0_d[20]) );
  CAOR2XL U343 ( .A(pushin), .B(q[21]), .C(n1431), .D(q0[21]), .Z(q0_d[21]) );
  CAOR2XL U342 ( .A(pushin), .B(q[22]), .C(n1432), .D(q0[22]), .Z(q0_d[22]) );
  CAOR2XL U341 ( .A(pushin), .B(q[23]), .C(n1432), .D(q0[23]), .Z(q0_d[23]) );
  CAOR2XL U332 ( .A(pushin), .B(h[0]), .C(n1430), .D(n419), .Z(h0_d[0]) );
  CAOR2XL U328 ( .A(pushin), .B(h[4]), .C(n1431), .D(n423), .Z(h0_d[4]) );
  CAOR2XL U327 ( .A(pushin), .B(h[5]), .C(n1431), .D(n424), .Z(h0_d[5]) );
  CAOR2XL U326 ( .A(pushin), .B(h[6]), .C(n1430), .D(n425), .Z(h0_d[6]) );
  CAOR2XL U329 ( .A(pushin), .B(h[3]), .C(n1432), .D(n422), .Z(h0_d[3]) );
  CAOR2XL U331 ( .A(pushin), .B(h[1]), .C(n1432), .D(n420), .Z(h0_d[1]) );
  CAOR2XL U330 ( .A(pushin), .B(h[2]), .C(n1431), .D(n421), .Z(h0_d[2]) );
  CND2XL \DP_OP_14_298_9081/U122  ( .A(\DP_OP_14_298_9081/n473 ), .B(
        \DP_OP_14_298_9081/n153 ), .Z(\DP_OP_14_298_9081/n16 ) );
  CND2XL \DP_OP_14_298_9081/U568  ( .A(\DP_OP_14_298_9081/n522 ), .B(
        \DP_OP_14_298_9081/n452 ), .Z(\DP_OP_14_298_9081/n65 ) );
  CND2XL \DP_OP_14_298_9081/U224  ( .A(\DP_OP_14_298_9081/n483 ), .B(
        \DP_OP_14_298_9081/n225 ), .Z(\DP_OP_14_298_9081/n26 ) );
  CND2XL \DP_OP_14_298_9081/U38  ( .A(\DP_OP_14_298_9081/n90 ), .B(
        \DP_OP_14_298_9081/n89 ), .Z(\DP_OP_14_298_9081/n8 ) );
  CND2XL \DP_OP_14_298_9081/U162  ( .A(\DP_OP_14_298_9081/n477 ), .B(
        \DP_OP_14_298_9081/n181 ), .Z(\DP_OP_14_298_9081/n20 ) );
  CND2XL \DP_OP_14_298_9081/U202  ( .A(\DP_OP_14_298_9081/n481 ), .B(
        \DP_OP_14_298_9081/n209 ), .Z(\DP_OP_14_298_9081/n24 ) );
  CND2XL \DP_OP_14_298_9081/U242  ( .A(\DP_OP_14_298_9081/n485 ), .B(
        \DP_OP_14_298_9081/n237 ), .Z(\DP_OP_14_298_9081/n28 ) );
  CND2XL \DP_OP_14_298_9081/U533  ( .A(\DP_OP_14_298_9081/n438 ), .B(
        \DP_OP_14_298_9081/n430 ), .Z(\DP_OP_14_298_9081/n428 ) );
  CND2XL \DP_OP_14_298_9081/U24  ( .A(\DP_OP_14_298_9081/n90 ), .B(n1190), .Z(
        \DP_OP_14_298_9081/n81 ) );
  CMX2XL U213 ( .A0(acc[20]), .A1(z[20]), .S(n201), .Z(n214) );
  CMX2XL U223 ( .A0(acc[10]), .A1(z[10]), .S(n201), .Z(n224) );
  CMX2XL U226 ( .A0(acc[7]), .A1(z[7]), .S(n201), .Z(n227) );
  CMX2XL U233 ( .A0(acc[0]), .A1(z[0]), .S(n201), .Z(n234) );
  CMX2XL U202 ( .A0(acc[31]), .A1(z[31]), .S(n201), .Z(n203) );
  CMX2XL U227 ( .A0(acc[6]), .A1(z[6]), .S(n201), .Z(n228) );
  CMX2XL U228 ( .A0(acc[5]), .A1(z[5]), .S(n201), .Z(n229) );
  CMX2XL U230 ( .A0(acc[3]), .A1(z[3]), .S(n201), .Z(n231) );
  CMX2XL U229 ( .A0(acc[4]), .A1(z[4]), .S(n201), .Z(n230) );
  CMX2XL U222 ( .A0(acc[11]), .A1(z[11]), .S(n201), .Z(n223) );
  CMX2XL U214 ( .A0(acc[19]), .A1(z[19]), .S(n201), .Z(n215) );
  CND2XL \DP_OP_14_298_9081/U264  ( .A(\DP_OP_14_298_9081/n487 ), .B(
        \DP_OP_14_298_9081/n253 ), .Z(\DP_OP_14_298_9081/n30 ) );
  CMX2XL U217 ( .A0(acc[16]), .A1(z[16]), .S(n201), .Z(n218) );
  CMX2XL U210 ( .A0(acc[23]), .A1(z[23]), .S(n201), .Z(n211) );
  CMX2XL U209 ( .A0(acc[24]), .A1(z[24]), .S(n201), .Z(n210) );
  CMX2XL U218 ( .A0(acc[15]), .A1(z[15]), .S(n201), .Z(n219) );
  CND2XL \DP_OP_14_298_9081/U12  ( .A(\DP_OP_14_298_9081/n463 ), .B(
        \DP_OP_14_298_9081/n73 ), .Z(\DP_OP_14_298_9081/n6 ) );
  CEOXL \DP_OP_14_298_9081/U578  ( .A(\DP_OP_14_298_9081/n461 ), .B(
        \DP_OP_14_298_9081/n67 ), .Z(\C1/DATA1_1 ) );
  CND2XL \DP_OP_14_298_9081/U318  ( .A(\DP_OP_14_298_9081/n493 ), .B(
        \DP_OP_14_298_9081/n289 ), .Z(\DP_OP_14_298_9081/n36 ) );
  COND1XL \DP_OP_14_298_9081/U465  ( .A(\DP_OP_14_298_9081/n385 ), .B(
        \DP_OP_14_298_9081/n406 ), .C(\DP_OP_14_298_9081/n386 ), .Z(
        \DP_OP_14_298_9081/n384 ) );
  CNR2XL \DP_OP_14_298_9081/U270  ( .A(\DP_OP_14_298_9081/n269 ), .B(
        \DP_OP_14_298_9081/n257 ), .Z(\DP_OP_14_298_9081/n255 ) );
  CND2XL \DP_OP_14_298_9081/U325  ( .A(\DP_OP_14_298_9081/n341 ), .B(
        \DP_OP_14_298_9081/n294 ), .Z(\DP_OP_14_298_9081/n292 ) );
  CND2XL \DP_OP_14_298_9081/U110  ( .A(\DP_OP_14_298_9081/n159 ), .B(
        \DP_OP_14_298_9081/n145 ), .Z(\DP_OP_14_298_9081/n143 ) );
  CND2XL \DP_OP_14_298_9081/U361  ( .A(\DP_OP_14_298_9081/n341 ), .B(
        \DP_OP_14_298_9081/n318 ), .Z(\DP_OP_14_298_9081/n316 ) );
  CEOXL \DP_OP_14_298_9081/U547  ( .A(\DP_OP_14_298_9081/n63 ), .B(
        \DP_OP_14_298_9081/n442 ), .Z(\C1/DATA1_5 ) );
  CNR2XL \DP_OP_14_298_9081/U86  ( .A(\DP_OP_14_298_9081/n4 ), .B(
        \DP_OP_14_298_9081/n127 ), .Z(\DP_OP_14_298_9081/n125 ) );
  CNR2XL \DP_OP_14_298_9081/U128  ( .A(\DP_OP_14_298_9081/n4 ), .B(
        \DP_OP_14_298_9081/n157 ), .Z(\DP_OP_14_298_9081/n155 ) );
  CNR2XL \DP_OP_14_298_9081/U108  ( .A(\DP_OP_14_298_9081/n4 ), .B(
        \DP_OP_14_298_9081/n143 ), .Z(\DP_OP_14_298_9081/n141 ) );
  CNR2XL \DP_OP_14_298_9081/U150  ( .A(\DP_OP_14_298_9081/n4 ), .B(
        \DP_OP_14_298_9081/n173 ), .Z(\DP_OP_14_298_9081/n171 ) );
  CNR2XL \DP_OP_14_298_9081/U66  ( .A(\DP_OP_14_298_9081/n4 ), .B(
        \DP_OP_14_298_9081/n113 ), .Z(\DP_OP_14_298_9081/n111 ) );
  CNR2XL \DP_OP_14_298_9081/U18  ( .A(\DP_OP_14_298_9081/n4 ), .B(
        \DP_OP_14_298_9081/n77 ), .Z(\DP_OP_14_298_9081/n75 ) );
  CNR2XL \DP_OP_14_298_9081/U190  ( .A(\DP_OP_14_298_9081/n213 ), .B(
        \DP_OP_14_298_9081/n201 ), .Z(\DP_OP_14_298_9081/n199 ) );
  CNR2XL \DP_OP_14_298_9081/U230  ( .A(\DP_OP_14_298_9081/n241 ), .B(
        \DP_OP_14_298_9081/n229 ), .Z(\DP_OP_14_298_9081/n227 ) );
  CEOXL \DP_OP_14_298_9081/U343  ( .A(\DP_OP_14_298_9081/n39 ), .B(
        \DP_OP_14_298_9081/n310 ), .Z(\C1/DATA1_29 ) );
  CAOR2XL U350 ( .A(pushin), .B(q[14]), .C(n1430), .D(q0[14]), .Z(q0_d[14]) );
  CAOR2XL U351 ( .A(pushin), .B(q[13]), .C(n1431), .D(q0[13]), .Z(q0_d[13]) );
  CND2XL \DP_OP_14_298_9081/U125  ( .A(acc[52]), .B(acc_a[52]), .Z(
        \DP_OP_14_298_9081/n153 ) );
  CND2XL \DP_OP_14_298_9081/U105  ( .A(acc[54]), .B(acc_a[54]), .Z(
        \DP_OP_14_298_9081/n139 ) );
  CAOR2XL U319 ( .A(pushin), .B(h[13]), .C(n1430), .D(h0[13]), .Z(h0_d[13]) );
  CAOR2XL U320 ( .A(pushin), .B(h[12]), .C(n1430), .D(h0[12]), .Z(h0_d[12]) );
  CAOR2XL U352 ( .A(pushin), .B(q[12]), .C(n1430), .D(q0[12]), .Z(q0_d[12]) );
  CAOR2XL U349 ( .A(pushin), .B(q[15]), .C(n1431), .D(q0[15]), .Z(q0_d[15]) );
  CAOR2XL U353 ( .A(pushin), .B(q[11]), .C(n1431), .D(q0[11]), .Z(q0_d[11]) );
  CND2XL \DP_OP_14_298_9081/U261  ( .A(acc[39]), .B(acc_a[39]), .Z(
        \DP_OP_14_298_9081/n250 ) );
  CAOR2XL U305 ( .A(pushin), .B(h[27]), .C(n1432), .D(h0[27]), .Z(h0_d[27]) );
  CND2XL \DP_OP_14_298_9081/U41  ( .A(acc[60]), .B(acc_a[60]), .Z(
        \DP_OP_14_298_9081/n89 ) );
  CAOR2XL U355 ( .A(pushin), .B(q[9]), .C(n1430), .D(q0[9]), .Z(q0_d[9]) );
  CAOR2XL U302 ( .A(pushin), .B(h[30]), .C(n1432), .D(h0[30]), .Z(h0_d[30]) );
  CND2XL \DP_OP_14_298_9081/U83  ( .A(n1087), .B(acc_a[56]), .Z(
        \DP_OP_14_298_9081/n123 ) );
  CAOR2XL U354 ( .A(pushin), .B(q[10]), .C(n1431), .D(q0[10]), .Z(q0_d[10]) );
  CND2XL \DP_OP_14_298_9081/U551  ( .A(\DP_OP_14_298_9081/n520 ), .B(
        \DP_OP_14_298_9081/n441 ), .Z(\DP_OP_14_298_9081/n63 ) );
  CND2XL \DP_OP_14_298_9081/U347  ( .A(\DP_OP_14_298_9081/n496 ), .B(
        \DP_OP_14_298_9081/n309 ), .Z(\DP_OP_14_298_9081/n39 ) );
  CND2XL \DP_OP_14_298_9081/U68  ( .A(\DP_OP_14_298_9081/n129 ), .B(
        \DP_OP_14_298_9081/n115 ), .Z(\DP_OP_14_298_9081/n113 ) );
  CNR2XL \DP_OP_14_298_9081/U22  ( .A(\DP_OP_14_298_9081/n101 ), .B(
        \DP_OP_14_298_9081/n81 ), .Z(\DP_OP_14_298_9081/n79 ) );
  CND2XL \DP_OP_14_298_9081/U46  ( .A(\DP_OP_14_298_9081/n129 ), .B(
        \DP_OP_14_298_9081/n99 ), .Z(\DP_OP_14_298_9081/n97 ) );
  CND2X1 \DP_OP_14_298_9081/U20  ( .A(\DP_OP_14_298_9081/n129 ), .B(
        \DP_OP_14_298_9081/n79 ), .Z(\DP_OP_14_298_9081/n77 ) );
  CND2XL \DP_OP_14_298_9081/U210  ( .A(\DP_OP_14_298_9081/n239 ), .B(
        \DP_OP_14_298_9081/n215 ), .Z(\DP_OP_14_298_9081/n213 ) );
  CANR1XL \DP_OP_14_298_9081/U481  ( .A(\DP_OP_14_298_9081/n395 ), .B(
        \DP_OP_14_298_9081/n404 ), .C(\DP_OP_14_298_9081/n396 ), .Z(
        \DP_OP_14_298_9081/n394 ) );
  CEOXL \DP_OP_14_298_9081/U480  ( .A(\DP_OP_14_298_9081/n55 ), .B(
        \DP_OP_14_298_9081/n399 ), .Z(\C1/DATA1_13 ) );
  CFD2XL \acc_reg[38]  ( .D(n158), .CP(clk), .CD(n199), .Q(n680), .QN(n679) );
  CFD4XL push2_reg ( .D(n428), .CP(clk), .SD(n199), .QN(n1417) );
  CFD4XL push1_reg ( .D(n430), .CP(clk), .SD(n199), .Q(n197), .QN(push1) );
  CFD4QXL push0_reg ( .D(n1431), .CP(clk), .SD(n199), .Q(n198) );
  CFD2QX1 \ho_2_reg[4]  ( .D(n432), .CP(clk), .CD(n199), .Q(ho_2[4]) );
  CFD3QX1 \acc_a_reg[23]  ( .D(n434), .CP(clk), .CD(n199), .SD(1'b1), .Q(
        acc_a[23]) );
  CFD2X4 \acc_reg[14]  ( .D(n182), .CP(clk), .CD(n199), .Q(n1095) );
  CENX1 \DP_OP_14_298_9081/U268  ( .A(\DP_OP_14_298_9081/n263 ), .B(
        \DP_OP_14_298_9081/n31 ), .Z(\C1/DATA1_37 ) );
  COND1XL \DP_OP_14_298_9081/U281  ( .A(\DP_OP_14_298_9081/n264 ), .B(
        \DP_OP_14_298_9081/n266 ), .C(\DP_OP_14_298_9081/n265 ), .Z(
        \DP_OP_14_298_9081/n263 ) );
  CND2X1 \DP_OP_14_298_9081/U276  ( .A(\DP_OP_14_298_9081/n488 ), .B(
        \DP_OP_14_298_9081/n262 ), .Z(\DP_OP_14_298_9081/n31 ) );
  CENX1 \DP_OP_14_298_9081/U308  ( .A(\DP_OP_14_298_9081/n287 ), .B(
        \DP_OP_14_298_9081/n35 ), .Z(\C1/DATA1_33 ) );
  COND1XL \DP_OP_14_298_9081/U317  ( .A(\DP_OP_14_298_9081/n288 ), .B(
        \DP_OP_14_298_9081/n290 ), .C(\DP_OP_14_298_9081/n289 ), .Z(
        \DP_OP_14_298_9081/n287 ) );
  CND2X1 \DP_OP_14_298_9081/U312  ( .A(\DP_OP_14_298_9081/n492 ), .B(
        \DP_OP_14_298_9081/n286 ), .Z(\DP_OP_14_298_9081/n35 ) );
  CFD2QX2 \acc_reg[25]  ( .D(n171), .CP(clk), .CD(n199), .Q(acc[25]) );
  CFD2QX2 \acc_reg[11]  ( .D(n185), .CP(clk), .CD(n199), .Q(acc[11]) );
  CFD2QX2 \acc_reg[31]  ( .D(n165), .CP(clk), .CD(n199), .Q(acc[31]) );
  CFD2QX2 \acc_reg[2]  ( .D(n194), .CP(clk), .CD(n199), .Q(acc[2]) );
  CFD2QX1 \acc_reg[48]  ( .D(n148), .CP(clk), .CD(n199), .Q(acc[48]) );
  CFD2QX2 \acc_reg[3]  ( .D(n193), .CP(clk), .CD(n199), .Q(acc[3]) );
  CEOXL \DP_OP_14_298_9081/U78  ( .A(\DP_OP_14_298_9081/n12 ), .B(
        \DP_OP_14_298_9081/n124 ), .Z(\C1/DATA1_56 ) );
  CND2XL \DP_OP_14_298_9081/U80  ( .A(\DP_OP_14_298_9081/n469 ), .B(
        \DP_OP_14_298_9081/n123 ), .Z(\DP_OP_14_298_9081/n12 ) );
  CENX1 \DP_OP_14_298_9081/U16  ( .A(\DP_OP_14_298_9081/n87 ), .B(
        \DP_OP_14_298_9081/n7 ), .Z(\C1/DATA1_61 ) );
  CND2X1 \DP_OP_14_298_9081/U28  ( .A(n1190), .B(\DP_OP_14_298_9081/n86 ), .Z(
        \DP_OP_14_298_9081/n7 ) );
  CEOXL \DP_OP_14_298_9081/U100  ( .A(\DP_OP_14_298_9081/n14 ), .B(
        \DP_OP_14_298_9081/n140 ), .Z(\C1/DATA1_54 ) );
  CND2XL \DP_OP_14_298_9081/U102  ( .A(\DP_OP_14_298_9081/n471 ), .B(
        \DP_OP_14_298_9081/n139 ), .Z(\DP_OP_14_298_9081/n14 ) );
  CFD2QX2 \acc_reg[42]  ( .D(n154), .CP(clk), .CD(n199), .Q(acc[42]) );
  CFD2X1 \acc_reg[45]  ( .D(n151), .CP(clk), .CD(n199), .Q(n309), .QN(n308) );
  CFD2QX2 \acc_reg[20]  ( .D(n176), .CP(clk), .CD(n199), .Q(acc[20]) );
  CFD2QX2 \acc_reg[54]  ( .D(n142), .CP(clk), .CD(n199), .Q(acc[54]) );
  CIVXL U366 ( .A(n816), .Z(n302) );
  COND1XL U367 ( .A(n1129), .B(n1513), .C(n1193), .Z(n1126) );
  CND2X1 U368 ( .A(n1333), .B(n1332), .Z(n1741) );
  CMXI2XL U369 ( .A0(acc[10]), .A1(acc[11]), .S(n435), .Z(n1540) );
  CNR2X4 U370 ( .A(n439), .B(n1026), .Z(n453) );
  CND2XL U371 ( .A(n777), .B(n1678), .Z(n822) );
  CMXI2XL U372 ( .A0(n1532), .A1(n1104), .S(n686), .Z(n1533) );
  CND3X1 U373 ( .A(n1707), .B(n1713), .C(n1705), .Z(n1648) );
  CIVXL U374 ( .A(n1415), .Z(n303) );
  CNR2X2 U375 ( .A(n304), .B(n305), .Z(n396) );
  CAN2X1 U376 ( .A(n777), .B(n1700), .Z(n304) );
  CAOR1X1 U377 ( .A(n1196), .B(\C1/DATA1_56 ), .C(n395), .Z(n305) );
  CND2X1 U378 ( .A(n348), .B(n349), .Z(n347) );
  CND3X2 U379 ( .A(n1003), .B(n1002), .C(n1784), .Z(n937) );
  CND2XL U380 ( .A(n838), .B(n1123), .Z(n306) );
  CND2XL U381 ( .A(n838), .B(n1123), .Z(n307) );
  CND2XL U382 ( .A(n838), .B(n1123), .Z(n1192) );
  CMXI2XL U383 ( .A0(n1516), .A1(n1517), .S(n1207), .Z(n1548) );
  CIVX2 U384 ( .A(n308), .Z(n310) );
  CMXI2XL U385 ( .A0(n1473), .A1(n642), .S(n1204), .Z(n416) );
  CMXI2XL U386 ( .A0(n641), .A1(n1473), .S(n544), .Z(n311) );
  CMXI2XL U387 ( .A0(n641), .A1(n1473), .S(n544), .Z(n1542) );
  CIVX1 U388 ( .A(n359), .Z(n887) );
  CND3X1 U389 ( .A(n338), .B(n1413), .C(n340), .Z(n337) );
  CNR2XL U390 ( .A(n1722), .B(n1911), .Z(n1721) );
  CANR1X1 U391 ( .A(n1422), .B(n1586), .C(n1411), .Z(n348) );
  CMXI2X1 U392 ( .A0(n1210), .A1(n351), .S(n367), .Z(n376) );
  CMXI2X2 U393 ( .A0(n1640), .A1(n1525), .S(n923), .Z(n1094) );
  CND3X1 U394 ( .A(n444), .B(n446), .C(n445), .Z(n312) );
  CMXI2X1 U395 ( .A0(n1526), .A1(n646), .S(n1422), .Z(n666) );
  CND3X1 U396 ( .A(n382), .B(n381), .C(n654), .Z(n313) );
  CND3X1 U397 ( .A(n654), .B(n381), .C(n382), .Z(n982) );
  CMXI2X1 U398 ( .A0(n1520), .A1(n341), .S(n542), .Z(n314) );
  CMXI2XL U399 ( .A0(n1520), .A1(n341), .S(n542), .Z(n343) );
  CNIVX4 U400 ( .A(ho_2[0]), .Z(n315) );
  CMXI2X1 U401 ( .A0(acc[48]), .A1(acc[49]), .S(n315), .Z(n1447) );
  CMXI2X1 U402 ( .A0(acc[50]), .A1(n1096), .S(n315), .Z(n1451) );
  CMXI2XL U403 ( .A0(n913), .A1(n914), .S(n315), .Z(n959) );
  CMXI2XL U404 ( .A0(acc[49]), .A1(acc[50]), .S(n315), .Z(n1472) );
  CMXI2X1 U405 ( .A0(n1096), .A1(acc[52]), .S(n315), .Z(n1471) );
  CMXI2XL U406 ( .A0(n916), .A1(acc[42]), .S(n315), .Z(n1470) );
  CMXI2XL U407 ( .A0(n917), .A1(acc[44]), .S(n315), .Z(n1469) );
  CMXI2XL U408 ( .A0(n309), .A1(acc[46]), .S(n315), .Z(n958) );
  CMXI2XL U409 ( .A0(n918), .A1(acc[48]), .S(n315), .Z(n1468) );
  CMXI2X1 U410 ( .A0(acc[53]), .A1(acc[54]), .S(n315), .Z(n1459) );
  CMXI2XL U411 ( .A0(acc[31]), .A1(n913), .S(n315), .Z(n1454) );
  CMXI2XL U412 ( .A0(n1438), .A1(n959), .S(n1420), .Z(n316) );
  CMXI2XL U413 ( .A0(n316), .A1(n1547), .S(n544), .Z(n321) );
  CND2IXL U414 ( .B(n316), .A(n1293), .Z(n961) );
  CND3X2 U415 ( .A(n880), .B(n317), .C(n1864), .Z(n874) );
  CENXL U416 ( .A(n317), .B(n1414), .Z(n1364) );
  CND2XL U417 ( .A(n1098), .B(n317), .Z(n1314) );
  CND2X2 U418 ( .A(n1113), .B(n1114), .Z(n317) );
  CMXI2XL U419 ( .A0(n1109), .A1(n1503), .S(n1203), .Z(n318) );
  CMXI2X1 U420 ( .A0(n318), .A1(n647), .S(n1427), .Z(n350) );
  CND2IXL U421 ( .B(n686), .A(n321), .Z(n320) );
  CANR1X1 U422 ( .A(n686), .B(n1624), .C(n1194), .Z(n319) );
  CND2X1 U423 ( .A(n319), .B(n320), .Z(n341) );
  CND2XL U424 ( .A(n350), .B(n1193), .Z(n649) );
  CMXI2X1 U425 ( .A0(n649), .A1(n1594), .S(n542), .Z(n1501) );
  CND3X1 U426 ( .A(n1107), .B(n1108), .C(n1426), .Z(n1861) );
  CND2X2 U427 ( .A(n1116), .B(n1103), .Z(n323) );
  CND2X2 U428 ( .A(n1861), .B(n1860), .Z(n322) );
  CND2X2 U429 ( .A(n322), .B(n323), .Z(n872) );
  CND2X2 U430 ( .A(n324), .B(n325), .Z(n1210) );
  CND2IX1 U431 ( .B(n544), .A(n1427), .Z(n328) );
  CND2X2 U432 ( .A(n1207), .B(n1427), .Z(n329) );
  CND2IXL U433 ( .B(ho_2[3]), .A(n1495), .Z(n330) );
  CND2X1 U434 ( .A(n330), .B(n331), .Z(n324) );
  CMXI2XL U435 ( .A0(n1454), .A1(n1463), .S(n547), .Z(n332) );
  CANR1XL U436 ( .A(ho_2[3]), .B(n332), .C(n1427), .Z(n331) );
  COND1XL U437 ( .A(n328), .B(n1608), .C(n1193), .Z(n327) );
  CNR2X1 U438 ( .A(n1497), .B(n329), .Z(n326) );
  CNR2X2 U439 ( .A(n326), .B(n327), .Z(n325) );
  CAN2XL U440 ( .A(n1712), .B(n1713), .Z(n333) );
  CND3XL U441 ( .A(n656), .B(n876), .C(n333), .Z(n1710) );
  CIVXL U442 ( .A(\DP_OP_14_298_9081/n138 ), .Z(\DP_OP_14_298_9081/n471 ) );
  CAOR2XL U443 ( .A(acc[54]), .B(n1416), .C(n1195), .D(acc_a[54]), .Z(n339) );
  CAN2XL U444 ( .A(n1711), .B(n1197), .Z(n340) );
  CIVXL U445 ( .A(n1710), .Z(n338) );
  CANR1XL U446 ( .A(n1196), .B(\C1/DATA1_54 ), .C(n339), .Z(n335) );
  CND2XL U447 ( .A(n777), .B(n1709), .Z(n336) );
  CND2XL U448 ( .A(n1710), .B(n1709), .Z(n334) );
  CND4X1 U449 ( .A(n337), .B(n334), .C(n336), .D(n335), .Z(n142) );
  CIVX2 U450 ( .A(n542), .Z(n342) );
  CND2X1 U451 ( .A(n341), .B(n342), .Z(n1107) );
  CND2IXL U452 ( .B(n1425), .A(n343), .Z(n346) );
  CND2X1 U453 ( .A(n314), .B(n1425), .Z(n1852) );
  CND2X1 U454 ( .A(n346), .B(n347), .Z(n344) );
  CND2X2 U455 ( .A(n344), .B(n1902), .Z(n345) );
  CIVXL U456 ( .A(n344), .Z(n1897) );
  CNR2X2 U457 ( .A(n357), .B(n345), .Z(n359) );
  CNR2X2 U458 ( .A(n357), .B(n345), .Z(n780) );
  CND2IXL U459 ( .B(n1422), .A(n1587), .Z(n349) );
  CND2IX1 U460 ( .B(n1429), .A(n350), .Z(n351) );
  CND2IX1 U461 ( .B(n543), .A(n351), .Z(n369) );
  CIVX2 U462 ( .A(n1421), .Z(n353) );
  CND3X1 U463 ( .A(n362), .B(n363), .C(n353), .Z(n354) );
  COND1X1 U464 ( .A(n353), .B(n1585), .C(n354), .Z(n375) );
  CANR1X1 U465 ( .A(n363), .B(n362), .C(n353), .Z(n352) );
  CANR1X1 U466 ( .A(n1030), .B(n1029), .C(n352), .Z(n1184) );
  CND2X2 U467 ( .A(n369), .B(n368), .Z(n355) );
  CND2X2 U468 ( .A(n355), .B(n1425), .Z(n379) );
  CNIVXL U469 ( .A(n355), .Z(n407) );
  CIVX2 U470 ( .A(n377), .Z(n356) );
  CND2X2 U471 ( .A(n356), .B(n370), .Z(n357) );
  CIVXL U472 ( .A(n356), .Z(n1906) );
  CIVX3 U473 ( .A(n380), .Z(n358) );
  CND2X1 U474 ( .A(n358), .B(n1182), .Z(n927) );
  CND2X2 U475 ( .A(n358), .B(n1182), .Z(n870) );
  CND2X1 U476 ( .A(n383), .B(n359), .Z(n360) );
  CAN2XL U477 ( .A(n780), .B(n1881), .Z(n1080) );
  CNR2X2 U478 ( .A(n655), .B(n360), .Z(n1098) );
  CNR2X2 U479 ( .A(n655), .B(n360), .Z(n657) );
  CIVX2 U480 ( .A(n871), .Z(n361) );
  CNR2X1 U481 ( .A(n361), .B(n874), .Z(n838) );
  CNR2X2 U482 ( .A(n361), .B(n874), .Z(n1146) );
  CMXI2XL U483 ( .A0(acc[11]), .A1(acc[12]), .S(n922), .Z(n1549) );
  CMXI2XL U484 ( .A0(n1549), .A1(n1554), .S(n1419), .Z(n1558) );
  CMXI2X1 U485 ( .A0(n1582), .A1(n1576), .S(n1419), .Z(n365) );
  CMXI2X1 U486 ( .A0(n365), .A1(n1558), .S(n545), .Z(n364) );
  CND2IX1 U487 ( .B(n686), .A(n364), .Z(n363) );
  CANR1X1 U488 ( .A(n686), .B(n1559), .C(n1429), .Z(n362) );
  CIVX2 U489 ( .A(n1421), .Z(n367) );
  CIVX2 U490 ( .A(n542), .Z(n366) );
  CANR2X1 U491 ( .A(n649), .B(n366), .C(n367), .D(n1594), .Z(n651) );
  CND2X1 U492 ( .A(n1210), .B(n543), .Z(n368) );
  CND2X2 U493 ( .A(n1894), .B(n1895), .Z(n370) );
  CND3X2 U494 ( .A(n372), .B(n371), .C(n1425), .Z(n1894) );
  CND2IX1 U495 ( .B(n373), .A(n1591), .Z(n372) );
  CIVX2 U496 ( .A(n543), .Z(n373) );
  CND2IX1 U497 ( .B(n374), .A(n1592), .Z(n371) );
  CIVX2 U498 ( .A(n1423), .Z(n374) );
  CMXI2X1 U499 ( .A0(n375), .A1(n376), .S(ho_2[4]), .Z(n377) );
  CND2X2 U500 ( .A(n1111), .B(n541), .Z(n378) );
  CND2X2 U501 ( .A(n379), .B(n378), .Z(n380) );
  CNR2X2 U502 ( .A(n1237), .B(n968), .Z(n382) );
  CNR2X2 U503 ( .A(n1240), .B(n1922), .Z(n381) );
  CNR2X1 U504 ( .A(n775), .B(n1145), .Z(n383) );
  COND1X1 U505 ( .A(\DP_OP_14_298_9081/n88 ), .B(\DP_OP_14_298_9081/n94 ), .C(
        \DP_OP_14_298_9081/n89 ), .Z(\DP_OP_14_298_9081/n87 ) );
  CANR2XL U506 ( .A(n1195), .B(acc_a[61]), .C(n1045), .D(n1416), .Z(n389) );
  CND2X1 U507 ( .A(\C1/DATA1_61 ), .B(n1196), .Z(n388) );
  CNR2IXL U508 ( .B(n1197), .A(n1675), .Z(n390) );
  CND2X1 U509 ( .A(n388), .B(n389), .Z(n387) );
  CIVXL U510 ( .A(n1674), .Z(n386) );
  CND2X1 U511 ( .A(n1414), .B(n390), .Z(n391) );
  CANR1XL U512 ( .A(n386), .B(n777), .C(n387), .Z(n385) );
  CND2IXL U513 ( .B(n391), .A(n1676), .Z(n384) );
  COND3XL U514 ( .A(n1676), .B(n1674), .C(n384), .D(n385), .Z(n135) );
  CIVXL U515 ( .A(\DP_OP_14_298_9081/n122 ), .Z(\DP_OP_14_298_9081/n469 ) );
  CAOR2XL U516 ( .A(n1087), .B(n1416), .C(n1195), .D(acc_a[56]), .Z(n395) );
  CIVXL U517 ( .A(n658), .Z(n394) );
  CND4XL U518 ( .A(n1414), .B(n658), .C(n1197), .D(n1701), .Z(n393) );
  CND2X1 U519 ( .A(n394), .B(n1700), .Z(n392) );
  CND3X1 U520 ( .A(n392), .B(n393), .C(n396), .Z(n140) );
  CND2X2 U521 ( .A(n1239), .B(n1238), .Z(n1240) );
  CNR2X1 U522 ( .A(n1240), .B(n1922), .Z(n397) );
  CND3X1 U523 ( .A(n1187), .B(n654), .C(n397), .Z(n655) );
  CNR2IXL U524 ( .B(\DP_OP_14_298_9081/n359 ), .A(\DP_OP_14_298_9081/n358 ), 
        .Z(n403) );
  CAOR2XL U525 ( .A(acc[20]), .B(n1416), .C(n1195), .D(acc_a[20]), .Z(n400) );
  CENX1 U526 ( .A(\DP_OP_14_298_9081/n360 ), .B(n403), .Z(\C1/DATA1_20 ) );
  CMXI2XL U527 ( .A0(n1078), .A1(n1857), .S(n1425), .Z(n401) );
  CND3XL U528 ( .A(n657), .B(n1056), .C(n1859), .Z(n402) );
  CANR1XL U529 ( .A(n1196), .B(\C1/DATA1_20 ), .C(n400), .Z(n399) );
  CENXL U530 ( .A(n402), .B(n401), .Z(n398) );
  COND1X1 U531 ( .A(n1911), .B(n398), .C(n399), .Z(n176) );
  CIVX8 U532 ( .A(n542), .Z(n1422) );
  CIVX2 U533 ( .A(n685), .Z(n534) );
  CIVX8 U534 ( .A(n543), .Z(n685) );
  CIVX3 U535 ( .A(n686), .Z(n464) );
  CIVX4 U536 ( .A(n1428), .Z(n1427) );
  COND3XL U537 ( .A(n1912), .B(n1911), .C(n557), .D(n1909), .Z(n192) );
  CNR2XL U538 ( .A(n1928), .B(n1922), .Z(n1918) );
  CENXL U539 ( .A(n1405), .B(n1918), .Z(n1919) );
  CENXL U540 ( .A(n1373), .B(n1374), .Z(n1368) );
  CND4X1 U541 ( .A(n1666), .B(n1667), .C(n1668), .D(n1665), .Z(n133) );
  CANR2X1 U542 ( .A(n1914), .B(n1927), .C(n1926), .D(\C1/DATA1_3 ), .Z(n1916)
         );
  COND1X1 U543 ( .A(n1416), .B(n1916), .C(n1915), .Z(n193) );
  CIVXL U544 ( .A(n1825), .Z(n1821) );
  COND1X1 U545 ( .A(n1416), .B(n1921), .C(n1920), .Z(n194) );
  COR2XL U546 ( .A(n1247), .B(n1661), .Z(n1005) );
  CND4XL U547 ( .A(n876), .B(n1796), .C(n1786), .D(n508), .Z(n404) );
  CND4XL U548 ( .A(n876), .B(n1796), .C(n1786), .D(n508), .Z(n877) );
  CIVX2 U549 ( .A(n1805), .Z(n834) );
  CND3X1 U550 ( .A(n667), .B(n1753), .C(n664), .Z(n405) );
  CNR2X2 U551 ( .A(n1693), .B(n1658), .Z(n1677) );
  CNR2XL U552 ( .A(n1751), .B(n1785), .Z(n1752) );
  COND3XL U553 ( .A(n1235), .B(n1911), .C(n1893), .D(n1892), .Z(n189) );
  CANR1X1 U554 ( .A(n1826), .B(n1825), .C(n1824), .Z(n1827) );
  CND4XL U555 ( .A(n442), .B(n441), .C(n678), .D(n1793), .Z(n406) );
  CND4XL U556 ( .A(n442), .B(n1793), .C(n678), .D(n441), .Z(n1792) );
  CND2IX2 U557 ( .B(n1412), .A(n1653), .Z(n1704) );
  CMXI2XL U558 ( .A0(acc[15]), .A1(acc[16]), .S(n1418), .Z(n1553) );
  CMXI2XL U559 ( .A0(acc[7]), .A1(acc[8]), .S(n1418), .Z(n1575) );
  CND2IX1 U560 ( .B(n541), .A(n1857), .Z(n1016) );
  CND2X1 U561 ( .A(n1857), .B(n541), .Z(n1895) );
  CNR2XL U562 ( .A(n853), .B(n1192), .Z(n847) );
  COND1X2 U563 ( .A(n1422), .B(n1627), .C(n971), .Z(n1655) );
  CMXI2XL U564 ( .A0(n1505), .A1(n1506), .S(n1207), .Z(n1062) );
  CMXI2XL U565 ( .A0(n1454), .A1(n1463), .S(n547), .Z(n408) );
  CIVXL U566 ( .A(n438), .Z(n1177) );
  CNR2X2 U567 ( .A(n1240), .B(n1922), .Z(n409) );
  CIVXL U568 ( .A(n1794), .Z(n410) );
  CIVXL U569 ( .A(n410), .Z(n411) );
  CNIVXL U570 ( .A(n1891), .Z(n412) );
  CIVXL U571 ( .A(n679), .Z(n681) );
  CND2XL U572 ( .A(n1224), .B(n1223), .Z(n413) );
  CND3X2 U573 ( .A(n453), .B(n945), .C(n1044), .Z(n1027) );
  CMX2GX2 U574 ( .GN(n1833), .A0(n466), .A1(n1831), .S(n1425), .Z(n945) );
  CMXI2X1 U575 ( .A0(n914), .A1(acc[34]), .S(n1418), .Z(n1463) );
  COR2X1 U576 ( .A(n1633), .B(n939), .Z(n507) );
  CIVXL U577 ( .A(n1640), .Z(n414) );
  CIVXL U578 ( .A(n414), .Z(n415) );
  CMXI2XL U579 ( .A0(n642), .A1(n1473), .S(n1424), .Z(n644) );
  CNIVX1 U580 ( .A(cmd1[1]), .Z(n417) );
  CNIVX3 U581 ( .A(cmd0[0]), .Z(n604) );
  CNIVX1 U582 ( .A(n604), .Z(n418) );
  CNIVXL U583 ( .A(h0[1]), .Z(n420) );
  CNIVXL U584 ( .A(h0[2]), .Z(n421) );
  CNIVXL U585 ( .A(h0[4]), .Z(n423) );
  CNIVXL U586 ( .A(h0[5]), .Z(n424) );
  CNIVXL U587 ( .A(h0[6]), .Z(n425) );
  CNIVXL U588 ( .A(h0[0]), .Z(n419) );
  CNIVXL U589 ( .A(h0[3]), .Z(n422) );
  CNIVX3 U590 ( .A(cmd0[1]), .Z(n635) );
  CNIVX1 U591 ( .A(n635), .Z(n426) );
  CNIVX3 U592 ( .A(h0_d_a[0]), .Z(n427) );
  CNIVX1 U593 ( .A(n429), .Z(n428) );
  CNIVX1 U594 ( .A(n197), .Z(n429) );
  CNIVX3 U595 ( .A(n198), .Z(n431) );
  CNIVX1 U596 ( .A(n431), .Z(n430) );
  CNIVX1 U597 ( .A(n433), .Z(n432) );
  CNIVX1 U598 ( .A(h0_d_a[4]), .Z(n433) );
  CNIVX1 U599 ( .A(n258), .Z(n434) );
  CNIVX4 U600 ( .A(ho_2[0]), .Z(n435) );
  CMXI2X1 U601 ( .A0(acc[58]), .A1(acc[59]), .S(n435), .Z(n770) );
  CMXI2XL U602 ( .A0(acc[3]), .A1(acc[4]), .S(n922), .Z(n1582) );
  CMXI2X1 U603 ( .A0(acc[20]), .A1(n1070), .S(n435), .Z(n1474) );
  CMXI2X1 U604 ( .A0(acc[52]), .A1(acc[53]), .S(n638), .Z(n639) );
  CMXI2X1 U605 ( .A0(acc[42]), .A1(n917), .S(n435), .Z(n1450) );
  CMXI2X1 U606 ( .A0(acc[46]), .A1(n918), .S(n435), .Z(n1448) );
  CMXI2X1 U607 ( .A0(acc[40]), .A1(n916), .S(n435), .Z(n1446) );
  CMXI2X1 U608 ( .A0(acc[60]), .A1(n1045), .S(n435), .Z(n1445) );
  CMXI2X1 U609 ( .A0(acc[30]), .A1(acc[31]), .S(n435), .Z(n1438) );
  CMXI2X1 U610 ( .A0(acc[24]), .A1(acc[25]), .S(n435), .Z(n1436) );
  CNR2IXL U611 ( .B(n1045), .A(n435), .Z(n898) );
  CND2IXL U612 ( .B(n1203), .A(n643), .Z(n436) );
  CND2IX1 U613 ( .B(n1280), .A(n436), .Z(n444) );
  CNR2X1 U614 ( .A(n1633), .B(n436), .Z(n1650) );
  CND3X2 U615 ( .A(n444), .B(n446), .C(n445), .Z(n437) );
  CMXI2X1 U616 ( .A0(n1210), .A1(n437), .S(n543), .Z(n448) );
  CMXI2X1 U617 ( .A0(n1210), .A1(n437), .S(n543), .Z(n1061) );
  CMXI2X1 U618 ( .A0(n312), .A1(n1642), .S(n1422), .Z(n1134) );
  CMXI2X1 U619 ( .A0(n312), .A1(n1642), .S(n1422), .Z(n1831) );
  CND2X2 U620 ( .A(n449), .B(n450), .Z(n438) );
  CND2X2 U621 ( .A(n1222), .B(n438), .Z(n439) );
  CND3X1 U622 ( .A(n1098), .B(n1183), .C(n438), .Z(n1400) );
  CNR2XL U623 ( .A(n439), .B(n1026), .Z(n1076) );
  CIVXL U624 ( .A(n439), .Z(n1849) );
  CND3X1 U625 ( .A(n453), .B(n945), .C(n1044), .Z(n440) );
  CNR2X2 U626 ( .A(n1410), .B(n440), .Z(n442) );
  CNR2X2 U627 ( .A(n1410), .B(n440), .Z(n912) );
  CNR2X2 U628 ( .A(n982), .B(n776), .Z(n441) );
  CND2XL U629 ( .A(n441), .B(n442), .Z(n1395) );
  CND3XL U630 ( .A(n442), .B(n441), .C(n1779), .Z(n1780) );
  CND3XL U631 ( .A(n441), .B(n458), .C(n442), .Z(n457) );
  CND3XL U632 ( .A(n442), .B(n441), .C(n1051), .Z(n1363) );
  CND3X1 U633 ( .A(n441), .B(n912), .C(n1793), .Z(n462) );
  CND3XL U634 ( .A(n656), .B(n441), .C(n912), .Z(n1736) );
  CND4XL U635 ( .A(n876), .B(n656), .C(n303), .D(n1662), .Z(n1666) );
  CIVXL U636 ( .A(n441), .Z(n1415) );
  CND3XL U637 ( .A(n1076), .B(n1851), .C(n441), .Z(n1841) );
  CND3XL U638 ( .A(n441), .B(n912), .C(n1796), .Z(n1797) );
  CND2XL U639 ( .A(n442), .B(n1098), .Z(n1377) );
  COND1X1 U640 ( .A(n1911), .B(n454), .C(n455), .Z(n163) );
  COND1X1 U641 ( .A(n1911), .B(n459), .C(n460), .Z(n159) );
  CMXI2XL U642 ( .A0(n1531), .A1(n1489), .S(n1424), .Z(n443) );
  CMXI2XL U643 ( .A0(n443), .A1(n772), .S(n686), .Z(n773) );
  CND2IX1 U644 ( .B(n686), .A(n1206), .Z(n447) );
  COAN1X1 U645 ( .A(n447), .B(n1502), .C(n1193), .Z(n445) );
  CND2IXL U646 ( .B(n1503), .A(n1293), .Z(n446) );
  CNR2IX1 U647 ( .B(n543), .A(n1525), .Z(n452) );
  CNR2X1 U648 ( .A(n1110), .B(n543), .Z(n451) );
  COND1X2 U649 ( .A(n451), .B(n452), .C(n1411), .Z(n450) );
  CND2IX1 U650 ( .B(n1411), .A(n448), .Z(n449) );
  CIVXL U651 ( .A(\DP_OP_14_298_9081/n285 ), .Z(\DP_OP_14_298_9081/n492 ) );
  CIVX1 U652 ( .A(n951), .Z(n458) );
  CAOR2XL U653 ( .A(n914), .B(n1416), .C(n1195), .D(acc_a[33]), .Z(n456) );
  CANR1XL U654 ( .A(n1196), .B(\C1/DATA1_33 ), .C(n456), .Z(n455) );
  CENXL U655 ( .A(n1803), .B(n457), .Z(n454) );
  CIVXL U656 ( .A(\DP_OP_14_298_9081/n261 ), .Z(\DP_OP_14_298_9081/n488 ) );
  CAOR2XL U657 ( .A(n944), .B(n1416), .C(n1195), .D(acc_a[37]), .Z(n461) );
  CANR1XL U658 ( .A(n1196), .B(\C1/DATA1_37 ), .C(n461), .Z(n460) );
  CEOXL U659 ( .A(n462), .B(n678), .Z(n459) );
  CMXI2X1 U660 ( .A0(n1515), .A1(n1484), .S(n1423), .Z(n934) );
  CIVDX4 U661 ( .A(n1193), .Z0(n1429) );
  CIVDX3 U662 ( .A(ho_2[6]), .Z0(n1193), .Z1(n1194) );
  CMXI2X1 U663 ( .A0(n867), .A1(n648), .S(n542), .Z(n650) );
  CMXI2X1 U664 ( .A0(n867), .A1(n1518), .S(n543), .Z(n868) );
  CMXI2X1 U665 ( .A0(n1528), .A1(n1118), .S(n464), .Z(n1117) );
  CNIVXL U666 ( .A(n1639), .Z(n465) );
  CMXI2XL U667 ( .A0(n1553), .A1(n1554), .S(n546), .Z(n1577) );
  CND2XL U668 ( .A(n1456), .B(n546), .Z(n1493) );
  CDLY1XL U669 ( .A(n1722), .Z(n1198) );
  COND1XL U670 ( .A(\DP_OP_14_298_9081/n405 ), .B(\DP_OP_14_298_9081/n426 ), 
        .C(\DP_OP_14_298_9081/n406 ), .Z(\DP_OP_14_298_9081/n404 ) );
  CND2X1 U671 ( .A(n1634), .B(n1422), .Z(n953) );
  COR2X1 U672 ( .A(n1426), .B(n1654), .Z(n1002) );
  CND2IX1 U673 ( .B(n1422), .A(n1598), .Z(n1131) );
  CANR1XL U674 ( .A(\DP_OP_14_298_9081/n353 ), .B(\DP_OP_14_298_9081/n361 ), 
        .C(\DP_OP_14_298_9081/n354 ), .Z(\DP_OP_14_298_9081/n352 ) );
  COND1XL U675 ( .A(\DP_OP_14_298_9081/n417 ), .B(\DP_OP_14_298_9081/n426 ), 
        .C(\DP_OP_14_298_9081/n418 ), .Z(\DP_OP_14_298_9081/n416 ) );
  COND1XL U676 ( .A(\DP_OP_14_298_9081/n245 ), .B(\DP_OP_14_298_9081/n270 ), 
        .C(\DP_OP_14_298_9081/n246 ), .Z(\DP_OP_14_298_9081/n240 ) );
  CANR1XL U677 ( .A(\DP_OP_14_298_9081/n513 ), .B(\DP_OP_14_298_9081/n404 ), 
        .C(\DP_OP_14_298_9081/n401 ), .Z(\DP_OP_14_298_9081/n399 ) );
  CND3XL U678 ( .A(n1774), .B(n1413), .C(n1071), .Z(n1775) );
  CAN2X1 U679 ( .A(n1926), .B(n1417), .Z(n1196) );
  CNR2IX1 U680 ( .B(cmd2[1]), .A(cmd2[0]), .Z(n1927) );
  CIVX2 U681 ( .A(n765), .Z(n1416) );
  CND3XL U682 ( .A(n684), .B(n1385), .C(n1383), .Z(n145) );
  CND2XL U683 ( .A(n1193), .B(n1427), .Z(n1031) );
  COND1XL U684 ( .A(n1193), .B(n1621), .C(n1423), .Z(n1034) );
  CMXI2XL U685 ( .A0(n1640), .A1(n1525), .S(n1423), .Z(n466) );
  CMXI2XL U686 ( .A0(n1111), .A1(n407), .S(n1425), .Z(n1859) );
  CND2XL U687 ( .A(\DP_OP_14_298_9081/n497 ), .B(\DP_OP_14_298_9081/n314 ), 
        .Z(n467) );
  CENXL U688 ( .A(\DP_OP_14_298_9081/n315 ), .B(n467), .Z(n468) );
  CND2X1 U689 ( .A(n1196), .B(n468), .Z(n1835) );
  CNR2IXL U690 ( .B(\DP_OP_14_298_9081/n351 ), .A(\DP_OP_14_298_9081/n350 ), 
        .Z(n469) );
  CENX1 U691 ( .A(\DP_OP_14_298_9081/n352 ), .B(n469), .Z(n470) );
  CND2X1 U692 ( .A(n1196), .B(n470), .Z(n902) );
  COND1XL U693 ( .A(\DP_OP_14_298_9081/n335 ), .B(\DP_OP_14_298_9081/n337 ), 
        .C(\DP_OP_14_298_9081/n336 ), .Z(n471) );
  CND2IXL U694 ( .B(\DP_OP_14_298_9081/n332 ), .A(\DP_OP_14_298_9081/n333 ), 
        .Z(n472) );
  CENX1 U695 ( .A(n471), .B(n472), .Z(\C1/DATA1_25 ) );
  CND2IX1 U696 ( .B(\DP_OP_14_298_9081/n264 ), .A(\DP_OP_14_298_9081/n265 ), 
        .Z(n473) );
  COND1XL U697 ( .A(n473), .B(\DP_OP_14_298_9081/n266 ), .C(n1196), .Z(n474)
         );
  CANR2XL U698 ( .A(acc[36]), .B(n1416), .C(acc_a[36]), .D(n1195), .Z(n475) );
  COND4CXL U699 ( .A(\DP_OP_14_298_9081/n266 ), .B(n473), .C(n474), .D(n475), 
        .Z(n1358) );
  CND2IXL U700 ( .B(\DP_OP_14_298_9081/n424 ), .A(\DP_OP_14_298_9081/n425 ), 
        .Z(n476) );
  COND1XL U701 ( .A(\DP_OP_14_298_9081/n426 ), .B(n476), .C(n1926), .Z(n477)
         );
  CANR1XL U702 ( .A(\DP_OP_14_298_9081/n426 ), .B(n476), .C(n477), .Z(n1200)
         );
  CMX2XL U703 ( .A0(n1570), .A1(n1547), .S(n545), .Z(n478) );
  CANR1X1 U704 ( .A(n686), .B(n1548), .C(n1429), .Z(n479) );
  COND1X1 U705 ( .A(n478), .B(n686), .C(n479), .Z(n1596) );
  COND1XL U706 ( .A(\DP_OP_14_298_9081/n369 ), .B(\DP_OP_14_298_9081/n371 ), 
        .C(\DP_OP_14_298_9081/n370 ), .Z(n480) );
  CND2IXL U707 ( .B(\DP_OP_14_298_9081/n366 ), .A(\DP_OP_14_298_9081/n367 ), 
        .Z(n481) );
  CENX1 U708 ( .A(n480), .B(n481), .Z(n803) );
  COND1XL U709 ( .A(\DP_OP_14_298_9081/n358 ), .B(\DP_OP_14_298_9081/n360 ), 
        .C(\DP_OP_14_298_9081/n359 ), .Z(n482) );
  CND2IXL U710 ( .B(\DP_OP_14_298_9081/n355 ), .A(\DP_OP_14_298_9081/n356 ), 
        .Z(n483) );
  CENX1 U711 ( .A(n482), .B(n483), .Z(n484) );
  CND2X1 U712 ( .A(n1196), .B(n484), .Z(n990) );
  CNR2IXL U713 ( .B(\DP_OP_14_298_9081/n422 ), .A(\DP_OP_14_298_9081/n421 ), 
        .Z(n485) );
  COND1XL U714 ( .A(\DP_OP_14_298_9081/n424 ), .B(\DP_OP_14_298_9081/n426 ), 
        .C(\DP_OP_14_298_9081/n425 ), .Z(n486) );
  COND1XL U715 ( .A(n485), .B(n486), .C(n1926), .Z(n487) );
  CANR1XL U716 ( .A(n485), .B(n486), .C(n487), .Z(n1199) );
  CND2IX1 U717 ( .B(\DP_OP_14_298_9081/n196 ), .A(\DP_OP_14_298_9081/n197 ), 
        .Z(n488) );
  COND1XL U718 ( .A(n488), .B(\DP_OP_14_298_9081/n198 ), .C(n1196), .Z(n489)
         );
  CANR2XL U719 ( .A(acc[46]), .B(n1416), .C(acc_a[46]), .D(n1195), .Z(n490) );
  COND4CXL U720 ( .A(\DP_OP_14_298_9081/n198 ), .B(n488), .C(n489), .D(n490), 
        .Z(n1299) );
  CANR2XL U721 ( .A(n1416), .B(acc[28]), .C(acc_a[28]), .D(n1195), .Z(n491) );
  CND2X1 U722 ( .A(n1835), .B(n491), .Z(n492) );
  CANR1XL U723 ( .A(n1837), .B(n1836), .C(n492), .Z(n1838) );
  CND2IX1 U724 ( .B(\DP_OP_14_298_9081/n327 ), .A(\DP_OP_14_298_9081/n328 ), 
        .Z(n493) );
  COND1XL U725 ( .A(n493), .B(\DP_OP_14_298_9081/n329 ), .C(n1196), .Z(n494)
         );
  CANR2XL U726 ( .A(acc[26]), .B(n1416), .C(acc_a[26]), .D(n1195), .Z(n495) );
  COND4CXL U727 ( .A(\DP_OP_14_298_9081/n329 ), .B(n493), .C(n494), .D(n495), 
        .Z(n1216) );
  CND3XL U728 ( .A(n1788), .B(n1106), .C(n1425), .Z(n1333) );
  CMXI2XL U729 ( .A0(n1638), .A1(n1637), .S(n1422), .Z(n496) );
  CAN2X1 U730 ( .A(n1425), .B(n496), .Z(n1731) );
  CNR2IXL U731 ( .B(\DP_OP_14_298_9081/n370 ), .A(\DP_OP_14_298_9081/n369 ), 
        .Z(n497) );
  CENX1 U732 ( .A(\DP_OP_14_298_9081/n371 ), .B(n497), .Z(n498) );
  CND2X1 U733 ( .A(n1196), .B(n498), .Z(n907) );
  CNR2IXL U734 ( .B(\DP_OP_14_298_9081/n336 ), .A(\DP_OP_14_298_9081/n335 ), 
        .Z(n499) );
  CENX1 U735 ( .A(\DP_OP_14_298_9081/n337 ), .B(n499), .Z(\C1/DATA1_24 ) );
  CND2XL U736 ( .A(\DP_OP_14_298_9081/n513 ), .B(\DP_OP_14_298_9081/n403 ), 
        .Z(n500) );
  CENX1 U737 ( .A(\DP_OP_14_298_9081/n404 ), .B(n500), .Z(n501) );
  CND2X1 U738 ( .A(n1926), .B(n501), .Z(n1337) );
  COND1XL U739 ( .A(\DP_OP_14_298_9081/n208 ), .B(\DP_OP_14_298_9081/n210 ), 
        .C(\DP_OP_14_298_9081/n209 ), .Z(n502) );
  CND2IXL U740 ( .B(\DP_OP_14_298_9081/n205 ), .A(\DP_OP_14_298_9081/n206 ), 
        .Z(n503) );
  CENXL U741 ( .A(n502), .B(n503), .Z(\C1/DATA1_45 ) );
  COND1XL U742 ( .A(\DP_OP_14_298_9081/n303 ), .B(\DP_OP_14_298_9081/n305 ), 
        .C(\DP_OP_14_298_9081/n304 ), .Z(n504) );
  CND2IXL U743 ( .B(\DP_OP_14_298_9081/n300 ), .A(\DP_OP_14_298_9081/n301 ), 
        .Z(n505) );
  CENX1 U744 ( .A(n504), .B(n505), .Z(\C1/DATA1_31 ) );
  CND2X1 U745 ( .A(n1848), .B(n1197), .Z(n506) );
  CNR2XL U746 ( .A(n1847), .B(n506), .Z(n1217) );
  CMXI2XL U747 ( .A0(n507), .A1(n1479), .S(n543), .Z(n1102) );
  COR2X1 U748 ( .A(n1412), .B(n954), .Z(n1735) );
  CNR2XL U749 ( .A(n1762), .B(n1765), .Z(n508) );
  CMX2XL U750 ( .A0(n1577), .A1(n1555), .S(n545), .Z(n509) );
  CANR1XL U751 ( .A(n686), .B(n962), .C(n1194), .Z(n510) );
  COND1XL U752 ( .A(n509), .B(n686), .C(n510), .Z(n963) );
  CANR2XL U753 ( .A(n1416), .B(acc[50]), .C(acc_a[50]), .D(n1195), .Z(n511) );
  CND2X1 U754 ( .A(n1403), .B(n511), .Z(n512) );
  CANR1XL U755 ( .A(n1728), .B(n1415), .C(n512), .Z(n1402) );
  CND2IXL U756 ( .B(n1147), .A(n1714), .Z(n826) );
  CIVX1 U757 ( .A(n1426), .Z(n513) );
  CNR2XL U758 ( .A(n1001), .B(n541), .Z(n514) );
  CANR1XL U759 ( .A(n1654), .B(n513), .C(n514), .Z(n949) );
  CND2X1 U760 ( .A(\DP_OP_14_298_9081/n509 ), .B(\DP_OP_14_298_9081/n381 ), 
        .Z(n515) );
  CND2XL U761 ( .A(n515), .B(\DP_OP_14_298_9081/n380 ), .Z(n516) );
  CND2IXL U762 ( .B(\DP_OP_14_298_9081/n374 ), .A(\DP_OP_14_298_9081/n375 ), 
        .Z(n517) );
  CENX1 U763 ( .A(n516), .B(n517), .Z(n518) );
  CND2X1 U764 ( .A(n1196), .B(n518), .Z(n985) );
  COND1XL U765 ( .A(\DP_OP_14_298_9081/n392 ), .B(\DP_OP_14_298_9081/n394 ), 
        .C(\DP_OP_14_298_9081/n393 ), .Z(n519) );
  CND2IXL U766 ( .B(\DP_OP_14_298_9081/n389 ), .A(\DP_OP_14_298_9081/n390 ), 
        .Z(n520) );
  CENX1 U767 ( .A(n519), .B(n520), .Z(\C1/DATA1_15 ) );
  COND1XL U768 ( .A(\DP_OP_14_298_9081/n350 ), .B(\DP_OP_14_298_9081/n352 ), 
        .C(\DP_OP_14_298_9081/n351 ), .Z(n521) );
  CND2IXL U769 ( .B(\DP_OP_14_298_9081/n347 ), .A(\DP_OP_14_298_9081/n348 ), 
        .Z(n522) );
  CENX1 U770 ( .A(n521), .B(n522), .Z(n1175) );
  CANR2XL U771 ( .A(acc[34]), .B(n1416), .C(acc_a[34]), .D(n1195), .Z(n523) );
  CND2IX1 U772 ( .B(\DP_OP_14_298_9081/n280 ), .A(\DP_OP_14_298_9081/n281 ), 
        .Z(n524) );
  COND1XL U773 ( .A(n524), .B(\DP_OP_14_298_9081/n282 ), .C(n1196), .Z(n525)
         );
  COND4CXL U774 ( .A(\DP_OP_14_298_9081/n282 ), .B(n524), .C(n525), .D(n523), 
        .Z(n1392) );
  CNR2IXL U775 ( .B(\DP_OP_14_298_9081/n304 ), .A(\DP_OP_14_298_9081/n303 ), 
        .Z(n526) );
  CENX1 U776 ( .A(\DP_OP_14_298_9081/n305 ), .B(n526), .Z(\C1/DATA1_30 ) );
  COND1XL U777 ( .A(\DP_OP_14_298_9081/n327 ), .B(\DP_OP_14_298_9081/n329 ), 
        .C(\DP_OP_14_298_9081/n328 ), .Z(n527) );
  CND2IXL U778 ( .B(\DP_OP_14_298_9081/n324 ), .A(\DP_OP_14_298_9081/n325 ), 
        .Z(n528) );
  CENX1 U779 ( .A(n527), .B(n528), .Z(\C1/DATA1_27 ) );
  CND2X1 U780 ( .A(\DP_OP_14_298_9081/n515 ), .B(\DP_OP_14_298_9081/n416 ), 
        .Z(n529) );
  CND2XL U781 ( .A(n529), .B(\DP_OP_14_298_9081/n415 ), .Z(n530) );
  CND2IXL U782 ( .B(\DP_OP_14_298_9081/n409 ), .A(\DP_OP_14_298_9081/n410 ), 
        .Z(n531) );
  CENX1 U783 ( .A(n530), .B(n531), .Z(\C1/DATA1_11 ) );
  CNR2IXL U784 ( .B(\DP_OP_14_298_9081/n436 ), .A(\DP_OP_14_298_9081/n435 ), 
        .Z(n532) );
  CENX1 U785 ( .A(\DP_OP_14_298_9081/n437 ), .B(n532), .Z(\C1/DATA1_6 ) );
  CNR2IXL U786 ( .B(\DP_OP_14_298_9081/n455 ), .A(\DP_OP_14_298_9081/n454 ), 
        .Z(n533) );
  CENX1 U787 ( .A(\DP_OP_14_298_9081/n456 ), .B(n533), .Z(\C1/DATA1_2 ) );
  CNR3XL U788 ( .A(n1552), .B(n1633), .C(n534), .Z(n1218) );
  CAOR1X1 U789 ( .A(n1275), .B(n1276), .C(n1423), .Z(n1150) );
  CND2IX1 U790 ( .B(\DP_OP_14_298_9081/n392 ), .A(\DP_OP_14_298_9081/n393 ), 
        .Z(n535) );
  COND1XL U791 ( .A(\DP_OP_14_298_9081/n394 ), .B(n535), .C(n1926), .Z(n536)
         );
  CANR1XL U792 ( .A(\DP_OP_14_298_9081/n394 ), .B(n535), .C(n536), .Z(n1868)
         );
  CAOR2X1 U793 ( .A(acc[19]), .B(n1416), .C(acc_a[19]), .D(n1195), .Z(n804) );
  CAOR1X1 U794 ( .A(n1196), .B(\C1/DATA1_52 ), .C(n1143), .Z(n537) );
  CANR1XL U795 ( .A(n777), .B(n1718), .C(n537), .Z(n1135) );
  COND1XL U796 ( .A(n1380), .B(n1192), .C(n1721), .Z(n1383) );
  CND2IX1 U797 ( .B(n1798), .A(n1796), .Z(n1357) );
  CAOR2X1 U798 ( .A(acc[15]), .B(n1416), .C(acc_a[15]), .D(n1195), .Z(n1366)
         );
  CAOR2X1 U799 ( .A(acc[23]), .B(n1416), .C(acc_a[23]), .D(n1195), .Z(n1176)
         );
  CAOR2X1 U800 ( .A(acc[24]), .B(n1416), .C(acc_a[24]), .D(n1195), .Z(n1398)
         );
  CIVX1 U801 ( .A(n1850), .Z(n538) );
  CND3XL U802 ( .A(n1851), .B(n1849), .C(n538), .Z(n1847) );
  CND2IX1 U803 ( .B(\DP_OP_14_298_9081/n432 ), .A(\DP_OP_14_298_9081/n433 ), 
        .Z(\DP_OP_14_298_9081/n61 ) );
  CND2IX1 U804 ( .B(\DP_OP_14_298_9081/n458 ), .A(\DP_OP_14_298_9081/n459 ), 
        .Z(\DP_OP_14_298_9081/n67 ) );
  COND1XL U805 ( .A(n1191), .B(n1725), .C(n1728), .Z(n539) );
  CND3XL U806 ( .A(n1401), .B(n1402), .C(n539), .Z(n146) );
  CIVDX1 U807 ( .A(n1411), .Z0(n540), .Z1(n541) );
  CIVDX1 U808 ( .A(n1911), .Z0(n1197) );
  CND2X2 U809 ( .A(n1927), .B(n1417), .Z(n1911) );
  CIVDX4 U810 ( .A(ho_2[2]), .Z0(n542), .Z1(n543) );
  CIVDX4 U811 ( .A(ho_2[3]), .Z0(n544), .Z1(n545) );
  CIVDX4 U812 ( .A(ho_2[1]), .Z0(n546), .Z1(n547) );
  CNIVX1 U813 ( .A(ho_2[4]), .Z(n1412) );
  CIVX4 U814 ( .A(n686), .Z(n1280) );
  CNIVXL U815 ( .A(n1887), .Z(n548) );
  CAN2X1 U816 ( .A(n1198), .B(n1197), .Z(n549) );
  CNR2X1 U817 ( .A(n1194), .B(n1427), .Z(n1035) );
  CNIVX1 U819 ( .A(n687), .Z(n552) );
  CNIVX1 U820 ( .A(n688), .Z(n553) );
  CNIVX1 U821 ( .A(n889), .Z(n554) );
  CNIVX1 U822 ( .A(n1899), .Z(n555) );
  CNIVX1 U823 ( .A(n1904), .Z(n556) );
  CNIVX1 U824 ( .A(n1910), .Z(n557) );
  CNIVX1 U825 ( .A(n250), .Z(n558) );
  CNIVX1 U826 ( .A(n251), .Z(n559) );
  CNIVX1 U827 ( .A(n252), .Z(n560) );
  CNIVX1 U828 ( .A(n253), .Z(n561) );
  CNIVX1 U829 ( .A(n254), .Z(n562) );
  CNIVX1 U830 ( .A(n255), .Z(n563) );
  CNIVX1 U831 ( .A(n256), .Z(n564) );
  CNIVX1 U832 ( .A(n257), .Z(n565) );
  CNIVX1 U833 ( .A(n259), .Z(n566) );
  CNIVX1 U834 ( .A(n260), .Z(n567) );
  CNIVX1 U835 ( .A(n261), .Z(n568) );
  CNIVX1 U836 ( .A(n262), .Z(n569) );
  CNIVX1 U837 ( .A(n263), .Z(n570) );
  CNIVX1 U838 ( .A(n264), .Z(n571) );
  CNIVX1 U839 ( .A(n265), .Z(n572) );
  CNIVX1 U840 ( .A(n266), .Z(n573) );
  CNIVX1 U841 ( .A(n267), .Z(n574) );
  CNIVX1 U842 ( .A(n268), .Z(n575) );
  CNIVX1 U843 ( .A(n269), .Z(n576) );
  CNIVX1 U844 ( .A(n270), .Z(n577) );
  CNIVX1 U845 ( .A(n271), .Z(n578) );
  CNIVX1 U846 ( .A(n272), .Z(n579) );
  CNIVX1 U847 ( .A(n273), .Z(n580) );
  CNIVX1 U848 ( .A(n274), .Z(n581) );
  CNIVX1 U849 ( .A(n275), .Z(n582) );
  CNIVX1 U850 ( .A(n276), .Z(n583) );
  CNIVX1 U851 ( .A(n277), .Z(n584) );
  CNIVX1 U852 ( .A(n278), .Z(n585) );
  CNIVX1 U853 ( .A(n279), .Z(n586) );
  CNIVX1 U854 ( .A(n280), .Z(n587) );
  CNIVX1 U855 ( .A(n281), .Z(n588) );
  CNIVX1 U856 ( .A(n282), .Z(n589) );
  CNIVX1 U857 ( .A(n283), .Z(n590) );
  CNIVX1 U858 ( .A(n284), .Z(n591) );
  CNIVX1 U859 ( .A(n285), .Z(n592) );
  CNIVX1 U860 ( .A(n286), .Z(n593) );
  CNIVX1 U861 ( .A(n288), .Z(n594) );
  CNIVX1 U862 ( .A(n289), .Z(n595) );
  CNIVX1 U863 ( .A(n290), .Z(n596) );
  CNIVX1 U864 ( .A(n292), .Z(n597) );
  CNIVX1 U865 ( .A(n293), .Z(n598) );
  CNIVX1 U866 ( .A(n294), .Z(n599) );
  CNIVX1 U867 ( .A(n700), .Z(n600) );
  CNIVX1 U868 ( .A(n702), .Z(n601) );
  CAN3X4 U869 ( .A(cmd2[0]), .B(cmd2[1]), .C(n765), .Z(_pushout_d) );
  CNIVX1 U870 ( .A(_pushout_d), .Z(n602) );
  CMX2X2 U871 ( .A0(n603), .A1(z[12]), .S(n201), .Z(n222) );
  CNIVX1 U872 ( .A(acc[12]), .Z(n603) );
  CNIVX1 U873 ( .A(n420), .Z(n605) );
  CNIVX1 U874 ( .A(n421), .Z(n606) );
  CNIVX1 U875 ( .A(n423), .Z(n607) );
  CNIVX1 U876 ( .A(n424), .Z(n608) );
  CNIVX1 U877 ( .A(n425), .Z(n609) );
  CNIVX1 U878 ( .A(n419), .Z(n610) );
  CNIVX1 U879 ( .A(n422), .Z(n611) );
  CMX2X2 U880 ( .A0(n612), .A1(z[1]), .S(n201), .Z(n233) );
  CNIVX1 U881 ( .A(acc[1]), .Z(n612) );
  CMX2X2 U882 ( .A0(n613), .A1(z[2]), .S(n201), .Z(n232) );
  CNIVX1 U883 ( .A(acc[2]), .Z(n613) );
  CNIVX1 U884 ( .A(n231), .Z(n614) );
  CNIVX1 U885 ( .A(n230), .Z(n615) );
  CNIVX1 U886 ( .A(n229), .Z(n616) );
  CNIVX1 U887 ( .A(n228), .Z(n617) );
  CNIVX1 U888 ( .A(n227), .Z(n618) );
  CMX2X2 U889 ( .A0(n763), .A1(z[8]), .S(n201), .Z(n226) );
  CMX2X2 U890 ( .A0(n761), .A1(z[9]), .S(n201), .Z(n225) );
  CNIVX1 U891 ( .A(n224), .Z(n619) );
  CNIVX1 U892 ( .A(n223), .Z(n620) );
  CMX2X2 U893 ( .A0(n766), .A1(z[13]), .S(n201), .Z(n221) );
  CMX2X2 U894 ( .A0(n1095), .A1(z[14]), .S(n201), .Z(n220) );
  CNIVX1 U895 ( .A(n219), .Z(n621) );
  CNIVX1 U896 ( .A(n218), .Z(n622) );
  CMX2X2 U897 ( .A0(n1069), .A1(z[17]), .S(n201), .Z(n217) );
  CMX2X2 U898 ( .A0(n1063), .A1(z[18]), .S(n201), .Z(n216) );
  CNIVX1 U899 ( .A(n215), .Z(n623) );
  CNIVX1 U900 ( .A(n214), .Z(n624) );
  CMX2X2 U901 ( .A0(n1070), .A1(z[21]), .S(n201), .Z(n213) );
  CMX2X2 U902 ( .A0(n1064), .A1(z[22]), .S(n201), .Z(n212) );
  CNIVX1 U903 ( .A(n211), .Z(n625) );
  CNIVX1 U904 ( .A(n210), .Z(n626) );
  CNIVX1 U905 ( .A(n209), .Z(n627) );
  CNIVX1 U906 ( .A(n208), .Z(n628) );
  CNIVX1 U907 ( .A(n207), .Z(n629) );
  CNIVX1 U908 ( .A(n206), .Z(n630) );
  CNIVX1 U909 ( .A(n205), .Z(n631) );
  CNIVX1 U910 ( .A(n204), .Z(n632) );
  CNIVX1 U911 ( .A(n203), .Z(n633) );
  CNIVX1 U912 ( .A(n234), .Z(n634) );
  CNIVX1 U913 ( .A(n760), .Z(n636) );
  CNIVX1 U914 ( .A(n768), .Z(n637) );
  CNIVX4 U915 ( .A(ho_2[0]), .Z(n638) );
  CMXI2XL U916 ( .A0(acc[34]), .A1(n915), .S(n638), .Z(n640) );
  CMXI2XL U917 ( .A0(n680), .A1(acc[39]), .S(n638), .Z(n864) );
  CMXI2XL U918 ( .A0(acc[9]), .A1(acc[10]), .S(n638), .Z(n1550) );
  CAN2XL U919 ( .A(n638), .B(n925), .Z(n899) );
  CANR1XL U920 ( .A(n638), .B(acc[0]), .C(n1419), .Z(n1037) );
  CMXI2XL U921 ( .A0(acc[25]), .A1(acc[26]), .S(n638), .Z(n1461) );
  CMXI2XL U922 ( .A0(acc[5]), .A1(acc[6]), .S(n638), .Z(n1576) );
  CMXI2XL U923 ( .A0(n1045), .A1(n925), .S(n638), .Z(n1457) );
  CMXI2X1 U924 ( .A0(n1087), .A1(n841), .S(n638), .Z(n1440) );
  CMXI2X1 U925 ( .A0(n841), .A1(acc[58]), .S(n638), .Z(n1465) );
  CMXI2X1 U926 ( .A0(acc[55]), .A1(n1087), .S(n638), .Z(n1208) );
  CMXI2X1 U927 ( .A0(n1070), .A1(n1064), .S(n638), .Z(n1453) );
  CMXI2X1 U928 ( .A0(n1451), .A1(n639), .S(n1420), .Z(n641) );
  CMXI2X1 U929 ( .A0(n1441), .A1(n639), .S(n546), .Z(n1505) );
  CMXI2X1 U930 ( .A0(n1444), .A1(n640), .S(n546), .Z(n642) );
  CMXI2X1 U931 ( .A0(n959), .A1(n640), .S(n1420), .Z(n1485) );
  CMXI2XL U932 ( .A0(n641), .A1(n1476), .S(n1424), .Z(n645) );
  COR2XL U933 ( .A(n1347), .B(n642), .Z(n1346) );
  COND1X1 U934 ( .A(n547), .B(n1464), .C(n897), .Z(n643) );
  CMXI2X1 U935 ( .A0(n1112), .A1(n643), .S(n1206), .Z(n647) );
  COR2X1 U936 ( .A(n1633), .B(n644), .Z(n648) );
  CMXI2X1 U937 ( .A0(n1273), .A1(n416), .S(n1427), .Z(n1272) );
  COR2X1 U938 ( .A(n1633), .B(n645), .Z(n646) );
  CANR1X1 U939 ( .A(n686), .B(n645), .C(n1194), .Z(n1232) );
  CMXI2X1 U940 ( .A0(n646), .A1(n1636), .S(n1422), .Z(n659) );
  CMXI2X1 U941 ( .A0(n646), .A1(n1636), .S(n1422), .Z(n910) );
  CMXI2XL U942 ( .A0(n1526), .A1(n646), .S(n1422), .Z(n1055) );
  COR2XL U943 ( .A(n1633), .B(n647), .Z(n1639) );
  CMXI2X1 U944 ( .A0(n1054), .A1(n648), .S(n1421), .Z(n1597) );
  CND2IXL U945 ( .B(n1411), .A(n650), .Z(n661) );
  CND2X1 U946 ( .A(n650), .B(n1411), .Z(n1860) );
  CMXI2X1 U947 ( .A0(n1184), .A1(n651), .S(n1411), .Z(n663) );
  CMXI2X1 U948 ( .A0(n1184), .A1(n651), .S(n1411), .Z(n1334) );
  CND2X1 U949 ( .A(n661), .B(n660), .Z(n652) );
  CND2X1 U950 ( .A(n1802), .B(n652), .Z(n662) );
  CNIVXL U951 ( .A(n652), .Z(n933) );
  CND2XL U952 ( .A(n413), .B(n652), .Z(n956) );
  CIVX2 U953 ( .A(n662), .Z(n653) );
  CND3X1 U954 ( .A(n653), .B(n941), .C(n1804), .Z(n1791) );
  CND4X1 U955 ( .A(n653), .B(n1161), .C(n932), .D(n1741), .Z(n1022) );
  CND4X1 U956 ( .A(n653), .B(n1161), .C(n932), .D(n1741), .Z(n818) );
  CNR2X2 U957 ( .A(n663), .B(n1917), .Z(n654) );
  CNR2X2 U958 ( .A(n1022), .B(n1018), .Z(n656) );
  CND3X1 U959 ( .A(n656), .B(n676), .C(n1101), .Z(n675) );
  CND4X1 U960 ( .A(n656), .B(n876), .C(n1101), .D(n1681), .Z(n1684) );
  CND4XL U961 ( .A(n1028), .B(n656), .C(n1101), .D(n1696), .Z(n1698) );
  CND2X1 U962 ( .A(n656), .B(n1101), .Z(n1379) );
  CND2XL U963 ( .A(n656), .B(n1381), .Z(n1380) );
  CND2IXL U964 ( .B(n1669), .A(n656), .Z(n1181) );
  CND3XL U965 ( .A(n657), .B(n1851), .C(n1849), .Z(n674) );
  CND2XL U966 ( .A(n657), .B(n1056), .Z(n806) );
  CND3XL U967 ( .A(n657), .B(n912), .C(n1763), .Z(n1764) );
  CND3XL U968 ( .A(n657), .B(n1856), .C(n1855), .Z(n904) );
  CND3XL U969 ( .A(n657), .B(n1863), .C(n1862), .Z(n909) );
  COND1X1 U970 ( .A(n1911), .B(n671), .C(n672), .Z(n171) );
  CNR2IX1 U971 ( .B(n1028), .A(n675), .Z(n658) );
  CND2IX1 U972 ( .B(n540), .A(n659), .Z(n660) );
  CNR2X1 U973 ( .A(n1649), .B(n1425), .Z(n670) );
  CAN2X1 U974 ( .A(n1017), .B(n1425), .Z(n669) );
  CANR2X1 U975 ( .A(n1094), .B(n669), .C(n670), .D(n1378), .Z(n668) );
  CMX2XL U976 ( .A0(n1660), .A1(n666), .S(n1426), .Z(n665) );
  CNR2X2 U977 ( .A(n1122), .B(n937), .Z(n664) );
  CNR2IX2 U978 ( .B(n665), .A(n668), .Z(n667) );
  CND3X2 U979 ( .A(n667), .B(n664), .C(n1753), .Z(n1018) );
  CAOR2XL U980 ( .A(acc[25]), .B(n1416), .C(n1195), .D(acc_a[25]), .Z(n673) );
  CANR1XL U981 ( .A(n1196), .B(\C1/DATA1_25 ), .C(n673), .Z(n672) );
  CENXL U982 ( .A(n674), .B(n1850), .Z(n671) );
  CIVXL U983 ( .A(n1704), .Z(n676) );
  CMXI2XL U984 ( .A0(n1497), .A1(n1608), .S(n545), .Z(n1632) );
  CNR3X1 U985 ( .A(n1791), .B(n1798), .C(n1795), .Z(n1793) );
  CNR3XL U986 ( .A(n1762), .B(n1791), .C(n1097), .Z(n1763) );
  CND2IXL U987 ( .B(n1791), .A(n1786), .Z(n1376) );
  CIVX2 U988 ( .A(n954), .Z(n677) );
  CND2X2 U989 ( .A(n952), .B(n953), .Z(n954) );
  CANR2X1 U990 ( .A(n1919), .B(n1927), .C(n1926), .D(\C1/DATA1_2 ), .Z(n1921)
         );
  CNIVXL U991 ( .A(n411), .Z(n678) );
  CND2IXL U992 ( .B(n1248), .A(n1703), .Z(n1011) );
  CANR1X2 U993 ( .A(n1293), .B(n1294), .C(n1194), .Z(n1289) );
  CND2X2 U994 ( .A(n1132), .B(n1133), .Z(n1085) );
  CMXI2X1 U995 ( .A0(n1502), .A1(n1504), .S(n1424), .Z(n1559) );
  CMXI2X1 U996 ( .A0(n1017), .A1(n1830), .S(n1426), .Z(n1833) );
  CND2X2 U997 ( .A(n1083), .B(n1084), .Z(n1079) );
  CAN2XL U998 ( .A(n1873), .B(n1187), .Z(n682) );
  CAN2XL U999 ( .A(n822), .B(n820), .Z(n683) );
  CAN2XL U1000 ( .A(n1384), .B(n1382), .Z(n684) );
  CND2XL U1001 ( .A(n777), .B(n1721), .Z(n1384) );
  CND2XL U1002 ( .A(n777), .B(n1703), .Z(n1012) );
  CNR2XL U1003 ( .A(n1252), .B(n1911), .Z(n1754) );
  CNR2XL U1004 ( .A(n1787), .B(n1911), .Z(n1375) );
  CND2IXL U1005 ( .B(n1848), .A(n1197), .Z(n1214) );
  CANR1XL U1006 ( .A(n1196), .B(n1175), .C(n1176), .Z(n1174) );
  CANR1XL U1007 ( .A(n1196), .B(n803), .C(n804), .Z(n802) );
  CNR2XL U1008 ( .A(n1715), .B(n1911), .Z(n1714) );
  CND2XL U1009 ( .A(n1081), .B(n1197), .Z(n1747) );
  CIVXL U1010 ( .A(n1679), .Z(n1672) );
  CNR2XL U1011 ( .A(n1671), .B(n1911), .Z(n1670) );
  CANR1X1 U1012 ( .A(n1422), .B(n1588), .C(n1411), .Z(n1139) );
  CND2XL U1013 ( .A(\C1/DATA1_4 ), .B(n1196), .Z(n1909) );
  CND2IXL U1014 ( .B(n1427), .A(n1320), .Z(n1319) );
  COND1XL U1015 ( .A(\DP_OP_14_298_9081/n131 ), .B(\DP_OP_14_298_9081/n158 ), 
        .C(\DP_OP_14_298_9081/n132 ), .Z(\DP_OP_14_298_9081/n130 ) );
  CIVXL U1016 ( .A(\DP_OP_14_298_9081/n320 ), .Z(\DP_OP_14_298_9081/n318 ) );
  CIVXL U1017 ( .A(\DP_OP_14_298_9081/n175 ), .Z(\DP_OP_14_298_9081/n173 ) );
  CANR2XL U1018 ( .A(n1195), .B(n701), .C(n603), .D(n1416), .Z(n1340) );
  CND2IXL U1019 ( .B(n686), .A(n545), .Z(n1347) );
  CIVXL U1020 ( .A(\DP_OP_14_298_9081/n259 ), .Z(\DP_OP_14_298_9081/n257 ) );
  CND2IXL U1021 ( .B(n686), .A(n545), .Z(n1351) );
  CIVXL U1022 ( .A(\DP_OP_14_298_9081/n203 ), .Z(\DP_OP_14_298_9081/n201 ) );
  CNR2X1 U1023 ( .A(n545), .B(n686), .Z(n1128) );
  CND2IXL U1024 ( .B(n686), .A(n1206), .Z(n1310) );
  CIVX2 U1025 ( .A(\DP_OP_14_298_9081/n89 ), .Z(\DP_OP_14_298_9081/n91 ) );
  CAN3X2 U1026 ( .A(n1434), .B(n1417), .C(n1433), .Z(n1195) );
  CIVXL U1027 ( .A(\DP_OP_14_298_9081/n88 ), .Z(\DP_OP_14_298_9081/n90 ) );
  CIVX1 U1028 ( .A(acc[63]), .Z(n1435) );
  CNR2X1 U1029 ( .A(n1095), .B(acc_a[14]), .Z(\DP_OP_14_298_9081/n392 ) );
  CND2XL U1030 ( .A(n1755), .B(n1754), .Z(n1758) );
  CENX1 U1031 ( .A(n1400), .B(n1399), .Z(n1396) );
  CND2IXL U1032 ( .B(n1214), .A(n1847), .Z(n1213) );
  CAN2XL U1033 ( .A(n1006), .B(n1004), .Z(n1009) );
  CIVXL U1034 ( .A(n1815), .Z(n1811) );
  CNR2XL U1035 ( .A(n1745), .B(n1744), .Z(n1746) );
  CNR2XL U1036 ( .A(n1376), .B(n793), .Z(n792) );
  CANR1XL U1037 ( .A(n1375), .B(n1376), .C(n786), .Z(n783) );
  CND2XL U1038 ( .A(n1393), .B(n1394), .Z(n1387) );
  CIVXL U1039 ( .A(n1391), .Z(n1393) );
  CIVXL U1040 ( .A(n1859), .Z(n805) );
  CNR2X1 U1041 ( .A(n950), .B(n956), .Z(n1796) );
  CIVXL U1042 ( .A(n1826), .Z(n1829) );
  CIVXL U1043 ( .A(n1375), .Z(n785) );
  CND2XL U1044 ( .A(n831), .B(n832), .Z(n830) );
  CIVXL U1045 ( .A(n1842), .Z(n1832) );
  CAN2X1 U1046 ( .A(n990), .B(n989), .Z(n849) );
  CIVXL U1047 ( .A(n1169), .Z(n1047) );
  CIVXL U1048 ( .A(n1214), .Z(n1215) );
  CIVXL U1049 ( .A(n1855), .Z(n991) );
  CND2XL U1050 ( .A(\C1/DATA1_63 ), .B(n1196), .Z(n1668) );
  CND2XL U1051 ( .A(n858), .B(n859), .Z(n857) );
  CAN2XL U1052 ( .A(n1686), .B(n1197), .Z(n840) );
  CND2XL U1053 ( .A(\C1/DATA1_53 ), .B(n1196), .Z(n831) );
  CIVX1 U1054 ( .A(n1862), .Z(n986) );
  CMXI2X1 U1055 ( .A0(n1053), .A1(n1788), .S(n540), .Z(n1798) );
  CAN2XL U1056 ( .A(n1072), .B(n1197), .Z(n1071) );
  CIVXL U1057 ( .A(n1837), .Z(n1840) );
  CND2XL U1058 ( .A(n1341), .B(n1417), .Z(n1339) );
  CNR2XL U1059 ( .A(n1735), .B(n1911), .Z(n1734) );
  CND2XL U1060 ( .A(n1371), .B(n1417), .Z(n1369) );
  CIVXL U1061 ( .A(n1694), .Z(n856) );
  CND2XL U1062 ( .A(\C1/DATA1_58 ), .B(n1196), .Z(n858) );
  CAN2XL U1063 ( .A(n1715), .B(n1197), .Z(n833) );
  CND2XL U1064 ( .A(\C1/DATA1_50 ), .B(n1196), .Z(n1403) );
  CIVXL U1065 ( .A(n1670), .Z(n1661) );
  CAN2XL U1066 ( .A(n1672), .B(n1675), .Z(n1180) );
  CND2XL U1067 ( .A(n1692), .B(n1685), .Z(n1658) );
  CMXI2X1 U1068 ( .A0(n1724), .A1(n929), .S(n1426), .Z(n1737) );
  CIVXL U1069 ( .A(n1868), .Z(n1872) );
  CAN2XL U1070 ( .A(n1699), .B(n1197), .Z(n1060) );
  CND2XL U1071 ( .A(n1823), .B(n1822), .Z(n1824) );
  CNR2XL U1072 ( .A(n1699), .B(n1911), .Z(n1697) );
  CAN2X1 U1073 ( .A(n985), .B(n984), .Z(n850) );
  CAN2X1 U1074 ( .A(n907), .B(n906), .Z(n896) );
  CIVXL U1075 ( .A(n1747), .Z(n1298) );
  CND2XL U1076 ( .A(n1685), .B(n1197), .Z(n1683) );
  CIVX1 U1077 ( .A(n1699), .Z(n1656) );
  CIVXL U1078 ( .A(n1876), .Z(n1880) );
  CAN2X1 U1079 ( .A(n902), .B(n901), .Z(n895) );
  CND2XL U1080 ( .A(n1337), .B(n1372), .Z(n1341) );
  CND2XL U1081 ( .A(\C1/DATA1_29 ), .B(n1196), .Z(n1823) );
  CNR2IXL U1082 ( .B(n1197), .A(n1081), .Z(n1300) );
  CNR2XL U1083 ( .A(n1711), .B(n1911), .Z(n1709) );
  CIVX1 U1084 ( .A(n1742), .Z(n1378) );
  CND2IX1 U1085 ( .B(n1425), .A(n1574), .Z(n1238) );
  CND2X1 U1086 ( .A(n1629), .B(n541), .Z(n1083) );
  CND2XL U1087 ( .A(n1675), .B(n1197), .Z(n1674) );
  CNR2XL U1088 ( .A(n1761), .B(n1911), .Z(n1760) );
  CND2XL U1089 ( .A(n1367), .B(n1372), .Z(n1371) );
  CND2XL U1090 ( .A(n1692), .B(n1197), .Z(n1694) );
  CND2XL U1091 ( .A(n1795), .B(n1197), .Z(n1359) );
  CIVXL U1092 ( .A(n1692), .Z(n1695) );
  CAN2XL U1093 ( .A(n1761), .B(n1197), .Z(n839) );
  CAN2XL U1094 ( .A(\C1/DATA1_11 ), .B(n1926), .Z(n892) );
  CAN2XL U1095 ( .A(\C1/DATA1_13 ), .B(n1926), .Z(n1876) );
  CNR2XL U1096 ( .A(n1795), .B(n1911), .Z(n1356) );
  CND2XL U1097 ( .A(n1660), .B(n1425), .Z(n1671) );
  CIVX1 U1098 ( .A(n1663), .Z(n1664) );
  CND2X1 U1099 ( .A(n976), .B(n977), .Z(n974) );
  CND2XL U1100 ( .A(\C1/DATA1_7 ), .B(n1196), .Z(n1892) );
  CANR1X1 U1101 ( .A(n1032), .B(n1033), .C(n1034), .Z(n1029) );
  CND2XL U1102 ( .A(\C1/DATA1_10 ), .B(n1926), .Z(n1367) );
  CIVXL U1103 ( .A(\DP_OP_14_298_9081/n4 ), .Z(\DP_OP_14_298_9081/n183 ) );
  CND2XL U1104 ( .A(\C1/DATA1_6 ), .B(n1196), .Z(n1898) );
  CND2XL U1105 ( .A(\C1/DATA1_5 ), .B(n1196), .Z(n1903) );
  CIVXL U1106 ( .A(\DP_OP_14_298_9081/n213 ), .Z(\DP_OP_14_298_9081/n211 ) );
  CIVXL U1107 ( .A(\DP_OP_14_298_9081/n269 ), .Z(\DP_OP_14_298_9081/n267 ) );
  CIVX1 U1108 ( .A(n1566), .Z(n1486) );
  CIVX1 U1109 ( .A(n1600), .Z(n1601) );
  CIVX1 U1110 ( .A(\DP_OP_14_298_9081/n101 ), .Z(\DP_OP_14_298_9081/n99 ) );
  CIVXL U1111 ( .A(\DP_OP_14_298_9081/n130 ), .Z(\DP_OP_14_298_9081/n128 ) );
  CND2IXL U1112 ( .B(n1427), .A(n1268), .Z(n1266) );
  CIVXL U1113 ( .A(\DP_OP_14_298_9081/n129 ), .Z(\DP_OP_14_298_9081/n127 ) );
  CIVXL U1114 ( .A(\DP_OP_14_298_9081/n158 ), .Z(\DP_OP_14_298_9081/n160 ) );
  CIVXL U1115 ( .A(\DP_OP_14_298_9081/n102 ), .Z(\DP_OP_14_298_9081/n100 ) );
  CIVXL U1116 ( .A(\DP_OP_14_298_9081/n157 ), .Z(\DP_OP_14_298_9081/n159 ) );
  CIVX1 U1117 ( .A(\DP_OP_14_298_9081/n217 ), .Z(\DP_OP_14_298_9081/n215 ) );
  CANR2XL U1118 ( .A(n1195), .B(acc_a[29]), .C(acc[29]), .D(n1416), .Z(n1822)
         );
  CIVXL U1119 ( .A(\DP_OP_14_298_9081/n288 ), .Z(\DP_OP_14_298_9081/n493 ) );
  CIVXL U1120 ( .A(\DP_OP_14_298_9081/n176 ), .Z(\DP_OP_14_298_9081/n174 ) );
  CANR2XL U1121 ( .A(n1195), .B(n691), .C(n612), .D(n1416), .Z(n1924) );
  CANR2XL U1122 ( .A(n1195), .B(n762), .C(n761), .D(n1416), .Z(n1884) );
  CANR2XL U1123 ( .A(n1195), .B(n769), .C(n1095), .D(n1416), .Z(n1869) );
  CANR2XL U1124 ( .A(n1195), .B(n767), .C(n766), .D(n1416), .Z(n1877) );
  CIVXL U1125 ( .A(n543), .Z(n1021) );
  CIVX2 U1126 ( .A(n543), .Z(n923) );
  CANR2XL U1127 ( .A(n1195), .B(n764), .C(n763), .D(n1416), .Z(n1889) );
  CANR2XL U1128 ( .A(n1195), .B(acc_a[22]), .C(n1064), .D(n1416), .Z(n901) );
  CIVXL U1129 ( .A(\DP_OP_14_298_9081/n260 ), .Z(\DP_OP_14_298_9081/n258 ) );
  CIVX1 U1130 ( .A(n1456), .Z(n1458) );
  CANR2XL U1131 ( .A(n1195), .B(acc_a[18]), .C(n1063), .D(n1416), .Z(n906) );
  CANR2XL U1132 ( .A(n1195), .B(acc_a[39]), .C(acc[39]), .D(n1416), .Z(n789)
         );
  CANR2XL U1133 ( .A(n1195), .B(n692), .C(n613), .D(n1416), .Z(n1920) );
  CANR2XL U1134 ( .A(n1195), .B(acc_a[53]), .C(acc[53]), .D(n1416), .Z(n832)
         );
  CANR2XL U1135 ( .A(n1195), .B(acc_a[63]), .C(acc[63]), .D(n1416), .Z(n1667)
         );
  CANR2XL U1136 ( .A(n1195), .B(acc_a[58]), .C(acc[58]), .D(n1416), .Z(n859)
         );
  CIVXL U1137 ( .A(\DP_OP_14_298_9081/n419 ), .Z(\DP_OP_14_298_9081/n417 ) );
  CIVXL U1138 ( .A(\DP_OP_14_298_9081/n204 ), .Z(\DP_OP_14_298_9081/n202 ) );
  CIVXL U1139 ( .A(\DP_OP_14_298_9081/n72 ), .Z(\DP_OP_14_298_9081/n463 ) );
  CANR2XL U1140 ( .A(n1195), .B(acc_a[17]), .C(n1069), .D(n1416), .Z(n984) );
  CIVXL U1141 ( .A(\DP_OP_14_298_9081/n231 ), .Z(\DP_OP_14_298_9081/n229 ) );
  CIVXL U1142 ( .A(\DP_OP_14_298_9081/n232 ), .Z(\DP_OP_14_298_9081/n230 ) );
  CIVXL U1143 ( .A(n1196), .Z(n787) );
  CANR2XL U1144 ( .A(n1195), .B(n693), .C(acc[3]), .D(n1416), .Z(n1915) );
  CANR2XL U1145 ( .A(n1195), .B(acc_a[21]), .C(n1070), .D(n1416), .Z(n989) );
  CND2XL U1146 ( .A(n542), .B(n1193), .Z(n1323) );
  CAN2XL U1147 ( .A(n1189), .B(\DP_OP_14_298_9081/n461 ), .Z(\C1/DATA1_0 ) );
  CIVX1 U1148 ( .A(\DP_OP_14_298_9081/n445 ), .Z(\DP_OP_14_298_9081/n521 ) );
  CIVXL U1149 ( .A(\DP_OP_14_298_9081/n446 ), .Z(\DP_OP_14_298_9081/n444 ) );
  CIVX1 U1150 ( .A(\DP_OP_14_298_9081/n403 ), .Z(\DP_OP_14_298_9081/n401 ) );
  CIVXL U1151 ( .A(\DP_OP_14_298_9081/n165 ), .Z(\DP_OP_14_298_9081/n474 ) );
  CIVX1 U1152 ( .A(\DP_OP_14_298_9081/n105 ), .Z(\DP_OP_14_298_9081/n466 ) );
  CIVXL U1153 ( .A(\DP_OP_14_298_9081/n180 ), .Z(\DP_OP_14_298_9081/n477 ) );
  CIVX1 U1154 ( .A(\DP_OP_14_298_9081/n313 ), .Z(\DP_OP_14_298_9081/n497 ) );
  CIVXL U1155 ( .A(\DP_OP_14_298_9081/n314 ), .Z(\DP_OP_14_298_9081/n312 ) );
  CIVXL U1156 ( .A(\DP_OP_14_298_9081/n308 ), .Z(\DP_OP_14_298_9081/n496 ) );
  CIVXL U1157 ( .A(\DP_OP_14_298_9081/n252 ), .Z(\DP_OP_14_298_9081/n487 ) );
  CIVXL U1158 ( .A(\DP_OP_14_298_9081/n119 ), .Z(\DP_OP_14_298_9081/n468 ) );
  CIVXL U1159 ( .A(\DP_OP_14_298_9081/n152 ), .Z(\DP_OP_14_298_9081/n473 ) );
  CND2IXL U1160 ( .B(\DP_OP_14_298_9081/n249 ), .A(\DP_OP_14_298_9081/n250 ), 
        .Z(n790) );
  CIVXL U1161 ( .A(\DP_OP_14_298_9081/n135 ), .Z(\DP_OP_14_298_9081/n470 ) );
  CIVXL U1162 ( .A(\DP_OP_14_298_9081/n236 ), .Z(\DP_OP_14_298_9081/n485 ) );
  CIVX1 U1163 ( .A(\DP_OP_14_298_9081/n402 ), .Z(\DP_OP_14_298_9081/n513 ) );
  CIVXL U1164 ( .A(\DP_OP_14_298_9081/n224 ), .Z(\DP_OP_14_298_9081/n483 ) );
  CIVXL U1165 ( .A(\DP_OP_14_298_9081/n208 ), .Z(\DP_OP_14_298_9081/n481 ) );
  CIVXL U1166 ( .A(\DP_OP_14_298_9081/n177 ), .Z(\DP_OP_14_298_9081/n476 ) );
  CIVX1 U1167 ( .A(\DP_OP_14_298_9081/n108 ), .Z(\DP_OP_14_298_9081/n467 ) );
  CIVXL U1168 ( .A(\DP_OP_14_298_9081/n86 ), .Z(\DP_OP_14_298_9081/n84 ) );
  CIVX1 U1169 ( .A(\DP_OP_14_298_9081/n149 ), .Z(\DP_OP_14_298_9081/n472 ) );
  CIVX1 U1170 ( .A(\DP_OP_14_298_9081/n233 ), .Z(\DP_OP_14_298_9081/n484 ) );
  CIVX1 U1171 ( .A(\DP_OP_14_298_9081/n379 ), .Z(\DP_OP_14_298_9081/n509 ) );
  CIVX1 U1172 ( .A(\DP_OP_14_298_9081/n414 ), .Z(\DP_OP_14_298_9081/n515 ) );
  CIVX1 U1173 ( .A(\DP_OP_14_298_9081/n221 ), .Z(\DP_OP_14_298_9081/n482 ) );
  CIVX1 U1174 ( .A(\DP_OP_14_298_9081/n168 ), .Z(\DP_OP_14_298_9081/n475 ) );
  CIVX1 U1175 ( .A(\DP_OP_14_298_9081/n193 ), .Z(\DP_OP_14_298_9081/n478 ) );
  CIVXL U1176 ( .A(\DP_OP_14_298_9081/n277 ), .Z(\DP_OP_14_298_9081/n490 ) );
  CIVX1 U1177 ( .A(n924), .Z(n926) );
  COR2XL U1178 ( .A(acc[63]), .B(acc_a[63]), .Z(n1188) );
  CIVX8 U1179 ( .A(n1428), .Z(n686) );
  COR2XL U1180 ( .A(acc[0]), .B(acc_a[0]), .Z(n1189) );
  CIVXL U1181 ( .A(n427), .Z(n931) );
  CNIVX1 U1182 ( .A(h0_d_a[5]), .Z(n687) );
  CNIVX1 U1183 ( .A(h0_d_a[6]), .Z(n688) );
  CANR2XL U1184 ( .A(n1195), .B(n699), .C(acc[11]), .D(n1416), .Z(n889) );
  CANR2XL U1185 ( .A(n1195), .B(n698), .C(acc[10]), .D(n1416), .Z(n1370) );
  CANR2XL U1186 ( .A(n1195), .B(n697), .C(acc[7]), .D(n1416), .Z(n1893) );
  CANR2XL U1187 ( .A(n1195), .B(n696), .C(acc[6]), .D(n1416), .Z(n1899) );
  CANR2XL U1188 ( .A(n1195), .B(n695), .C(acc[5]), .D(n1416), .Z(n1904) );
  CANR2XL U1189 ( .A(n1195), .B(n694), .C(acc[4]), .D(n1416), .Z(n1910) );
  CNIVX1 U1190 ( .A(n196), .Z(n689) );
  CANR2XL U1191 ( .A(n1195), .B(n690), .C(acc[0]), .D(n1416), .Z(n1931) );
  CNIVX1 U1192 ( .A(acc_a[0]), .Z(n690) );
  CNIVX1 U1193 ( .A(acc_a[1]), .Z(n691) );
  CNIVX1 U1194 ( .A(acc_a[2]), .Z(n692) );
  CNIVX1 U1195 ( .A(acc_a[3]), .Z(n693) );
  CNIVX1 U1196 ( .A(acc_a[4]), .Z(n694) );
  CNIVX1 U1197 ( .A(acc_a[5]), .Z(n695) );
  CNIVX1 U1198 ( .A(acc_a[6]), .Z(n696) );
  CNIVX1 U1199 ( .A(acc_a[7]), .Z(n697) );
  CNIVX1 U1200 ( .A(acc_a[10]), .Z(n698) );
  CNIVX1 U1201 ( .A(acc_a[11]), .Z(n699) );
  CNIVX1 U1202 ( .A(cmd1[0]), .Z(n700) );
  CNIVX1 U1203 ( .A(acc_a[12]), .Z(n701) );
  CNIVX1 U1204 ( .A(h0_d_a[3]), .Z(n702) );
  CNIVX1 U1205 ( .A(q0_d[0]), .Z(n703) );
  CNIVX1 U1206 ( .A(h0_d[7]), .Z(n704) );
  CNIVX1 U1207 ( .A(h0_d[8]), .Z(n705) );
  CNIVX1 U1208 ( .A(h0_d[9]), .Z(n706) );
  CNIVX1 U1209 ( .A(h0_d[10]), .Z(n707) );
  CNIVX1 U1210 ( .A(h0_d[11]), .Z(n708) );
  CNIVX1 U1211 ( .A(h0_d[12]), .Z(n709) );
  CNIVX1 U1212 ( .A(h0_d[13]), .Z(n710) );
  CNIVX1 U1213 ( .A(h0_d[14]), .Z(n711) );
  CNIVX1 U1214 ( .A(h0_d[15]), .Z(n712) );
  CNIVX1 U1215 ( .A(h0_d[16]), .Z(n713) );
  CNIVX1 U1216 ( .A(h0_d[17]), .Z(n714) );
  CNIVX1 U1217 ( .A(h0_d[18]), .Z(n715) );
  CNIVX1 U1218 ( .A(h0_d[19]), .Z(n716) );
  CNIVX1 U1219 ( .A(h0_d[20]), .Z(n717) );
  CNIVX1 U1220 ( .A(h0_d[21]), .Z(n718) );
  CNIVX1 U1221 ( .A(h0_d[22]), .Z(n719) );
  CNIVX1 U1222 ( .A(h0_d[23]), .Z(n720) );
  CNIVX1 U1223 ( .A(h0_d[24]), .Z(n721) );
  CNIVX1 U1224 ( .A(h0_d[25]), .Z(n722) );
  CNIVX1 U1225 ( .A(h0_d[26]), .Z(n723) );
  CNIVX1 U1226 ( .A(h0_d[27]), .Z(n724) );
  CNIVX1 U1227 ( .A(h0_d[28]), .Z(n725) );
  CNIVX1 U1228 ( .A(h0_d[29]), .Z(n726) );
  CNIVX1 U1229 ( .A(h0_d[30]), .Z(n727) );
  CNIVX1 U1230 ( .A(h0_d[31]), .Z(n728) );
  CNIVX1 U1231 ( .A(q0_d[1]), .Z(n729) );
  CNIVX1 U1232 ( .A(q0_d[2]), .Z(n730) );
  CNIVX1 U1233 ( .A(q0_d[3]), .Z(n731) );
  CNIVX1 U1234 ( .A(q0_d[4]), .Z(n732) );
  CNIVX1 U1235 ( .A(q0_d[5]), .Z(n733) );
  CNIVX1 U1236 ( .A(q0_d[6]), .Z(n734) );
  CNIVX1 U1237 ( .A(q0_d[7]), .Z(n735) );
  CNIVX1 U1238 ( .A(q0_d[8]), .Z(n736) );
  CNIVX1 U1239 ( .A(q0_d[9]), .Z(n737) );
  CNIVX1 U1240 ( .A(q0_d[10]), .Z(n738) );
  CNIVX1 U1241 ( .A(q0_d[11]), .Z(n739) );
  CNIVX1 U1242 ( .A(q0_d[12]), .Z(n740) );
  CNIVX1 U1243 ( .A(q0_d[13]), .Z(n741) );
  CNIVX1 U1244 ( .A(q0_d[14]), .Z(n742) );
  CNIVX1 U1245 ( .A(q0_d[15]), .Z(n743) );
  CNIVX1 U1246 ( .A(q0_d[16]), .Z(n744) );
  CNIVX1 U1247 ( .A(q0_d[17]), .Z(n745) );
  CNIVX1 U1248 ( .A(q0_d[18]), .Z(n746) );
  CNIVX1 U1249 ( .A(q0_d[19]), .Z(n747) );
  CNIVX1 U1250 ( .A(q0_d[20]), .Z(n748) );
  CNIVX1 U1251 ( .A(q0_d[21]), .Z(n749) );
  CNIVX1 U1252 ( .A(q0_d[22]), .Z(n750) );
  CNIVX1 U1253 ( .A(q0_d[23]), .Z(n751) );
  CNIVX1 U1254 ( .A(q0_d[24]), .Z(n752) );
  CNIVX1 U1255 ( .A(q0_d[25]), .Z(n753) );
  CNIVX1 U1256 ( .A(q0_d[26]), .Z(n754) );
  CNIVX1 U1257 ( .A(q0_d[27]), .Z(n755) );
  CNIVX1 U1258 ( .A(q0_d[28]), .Z(n756) );
  CNIVX1 U1259 ( .A(q0_d[29]), .Z(n757) );
  CNIVX1 U1260 ( .A(q0_d[30]), .Z(n758) );
  CNIVX1 U1261 ( .A(q0_d[31]), .Z(n759) );
  CNIVX1 U1262 ( .A(h0_d_a[1]), .Z(n760) );
  CNIVX1 U1263 ( .A(acc[9]), .Z(n761) );
  CNIVX1 U1264 ( .A(acc_a[9]), .Z(n762) );
  CNIVX1 U1265 ( .A(acc[8]), .Z(n763) );
  CNIVX1 U1266 ( .A(acc_a[8]), .Z(n764) );
  CNIVX1 U1267 ( .A(n1417), .Z(n765) );
  CNIVX1 U1268 ( .A(acc[13]), .Z(n766) );
  CNIVX1 U1269 ( .A(acc_a[13]), .Z(n767) );
  CNIVX1 U1270 ( .A(h0_d_a[2]), .Z(n768) );
  CNIVX1 U1271 ( .A(acc_a[14]), .Z(n769) );
  CIVX8 U1272 ( .A(rst), .Z(n199) );
  CMXI2X1 U1273 ( .A0(n1440), .A1(n770), .S(n1420), .Z(n771) );
  CMXI2X1 U1274 ( .A0(n770), .A1(n1445), .S(n1420), .Z(n1476) );
  CMXI2XL U1275 ( .A0(n1490), .A1(n771), .S(n1206), .Z(n772) );
  CND2IXL U1276 ( .B(n1203), .A(n771), .Z(n1605) );
  COR2XL U1277 ( .A(n1633), .B(n772), .Z(n1631) );
  CND2IXL U1278 ( .B(n1194), .A(n773), .Z(n779) );
  CND2IXL U1279 ( .B(n1194), .A(n773), .Z(n919) );
  CMX2X2 U1280 ( .A0(n778), .A1(n1830), .S(n1411), .Z(n774) );
  CND2X2 U1281 ( .A(n774), .B(n1085), .Z(n775) );
  CIVXL U1282 ( .A(n774), .Z(n1342) );
  CNR2X2 U1283 ( .A(n775), .B(n1145), .Z(n781) );
  CIVXL U1284 ( .A(n775), .Z(n1873) );
  CND2X2 U1285 ( .A(n781), .B(n780), .Z(n776) );
  CNR2X2 U1286 ( .A(n313), .B(n776), .Z(n969) );
  CIVX2 U1287 ( .A(n969), .Z(n777) );
  CND2XL U1288 ( .A(n777), .B(n1732), .Z(n796) );
  CANR1XL U1289 ( .A(n1714), .B(n777), .C(n830), .Z(n827) );
  CANR1XL U1290 ( .A(n856), .B(n777), .C(n857), .Z(n855) );
  CND2XL U1291 ( .A(n777), .B(n1760), .Z(n883) );
  CND2XL U1292 ( .A(n777), .B(n1814), .Z(n1817) );
  CND2XL U1293 ( .A(n777), .B(n1754), .Z(n1757) );
  CND2XL U1294 ( .A(n777), .B(n1697), .Z(n1154) );
  CND2XL U1295 ( .A(n777), .B(n1670), .Z(n1006) );
  CANR1XL U1296 ( .A(n1298), .B(n777), .C(n1299), .Z(n1297) );
  CANR1XL U1297 ( .A(n1215), .B(n777), .C(n1216), .Z(n1212) );
  CMXI2X1 U1298 ( .A0(n1593), .A1(n779), .S(ho_2[2]), .Z(n778) );
  CND2IX1 U1299 ( .B(n1911), .A(n1787), .Z(n793) );
  CND2IXL U1300 ( .B(n785), .A(n1377), .Z(n784) );
  CND3XL U1301 ( .A(n782), .B(n784), .C(n783), .Z(n157) );
  COAN1XL U1302 ( .A(\DP_OP_14_298_9081/n252 ), .B(\DP_OP_14_298_9081/n254 ), 
        .C(\DP_OP_14_298_9081/n253 ), .Z(n791) );
  CENXL U1303 ( .A(n790), .B(n791), .Z(n788) );
  CND2IXL U1304 ( .B(n1377), .A(n792), .Z(n782) );
  COND1XL U1305 ( .A(n787), .B(n788), .C(n789), .Z(n786) );
  CAOR2XL U1306 ( .A(acc[49]), .B(n1416), .C(n1195), .D(acc_a[49]), .Z(n799)
         );
  CIVXL U1307 ( .A(n1158), .Z(n798) );
  CANR1XL U1308 ( .A(n1196), .B(\C1/DATA1_49 ), .C(n799), .Z(n794) );
  CND2X1 U1309 ( .A(n798), .B(n1732), .Z(n795) );
  CND4XL U1310 ( .A(n1158), .B(n1413), .C(n1197), .D(n1733), .Z(n797) );
  CAN2X1 U1311 ( .A(n796), .B(n794), .Z(n800) );
  CND3X1 U1312 ( .A(n800), .B(n797), .C(n795), .Z(n147) );
  CENXL U1313 ( .A(n806), .B(n805), .Z(n801) );
  COND1X1 U1314 ( .A(n1911), .B(n801), .C(n802), .Z(n177) );
  CND2IXL U1315 ( .B(n1737), .A(n846), .Z(n807) );
  COND1XL U1316 ( .A(n807), .B(n1191), .C(n1734), .Z(n809) );
  CNR2XL U1317 ( .A(n306), .B(n807), .Z(n813) );
  CND4XL U1318 ( .A(n811), .B(n808), .C(n810), .D(n809), .Z(n148) );
  CAOR2XL U1319 ( .A(acc[48]), .B(n1416), .C(n1195), .D(acc_a[48]), .Z(n812)
         );
  CND4XL U1320 ( .A(n813), .B(n1414), .C(n1197), .D(n1735), .Z(n811) );
  CND2XL U1321 ( .A(n1415), .B(n1734), .Z(n810) );
  CANR1XL U1322 ( .A(n1196), .B(\C1/DATA1_48 ), .C(n812), .Z(n808) );
  CMX2X1 U1323 ( .A0(n1271), .A1(n1587), .S(n1422), .Z(n1270) );
  CIVX2 U1324 ( .A(n1075), .Z(n1628) );
  CND2X2 U1325 ( .A(n1887), .B(n1236), .Z(n1237) );
  CND2IX1 U1326 ( .B(n814), .A(n1891), .Z(n1886) );
  CIVXL U1327 ( .A(n1236), .Z(n814) );
  COND4CX1 U1328 ( .A(n1927), .B(n1888), .C(n1200), .D(n765), .Z(n1890) );
  CND2IXL U1329 ( .B(n815), .A(n846), .Z(n819) );
  CIVXL U1330 ( .A(n1712), .Z(n815) );
  CND2X2 U1331 ( .A(n1794), .B(n845), .Z(n816) );
  CIVXL U1332 ( .A(n816), .Z(n817) );
  CIVX2 U1333 ( .A(n816), .Z(n932) );
  CND3X1 U1334 ( .A(n823), .B(n683), .C(n821), .Z(n136) );
  CNR2X2 U1335 ( .A(n405), .B(n818), .Z(n846) );
  CNR2X1 U1336 ( .A(n1191), .B(n819), .Z(n1147) );
  CAOR2XL U1337 ( .A(acc[60]), .B(n1416), .C(n1195), .D(acc_a[60]), .Z(n825)
         );
  CANR1XL U1338 ( .A(n1196), .B(\C1/DATA1_60 ), .C(n825), .Z(n820) );
  CIVXL U1339 ( .A(n1680), .Z(n824) );
  CND4XL U1340 ( .A(n1680), .B(n1414), .C(n1197), .D(n1679), .Z(n823) );
  CND2X1 U1341 ( .A(n824), .B(n1678), .Z(n821) );
  CENXL U1342 ( .A(\DP_OP_14_298_9081/n151 ), .B(\DP_OP_14_298_9081/n15 ), .Z(
        \C1/DATA1_53 ) );
  CND2XL U1343 ( .A(n1414), .B(n833), .Z(n829) );
  CND2IXL U1344 ( .B(n829), .A(n1147), .Z(n828) );
  CND3XL U1345 ( .A(n826), .B(n828), .C(n827), .Z(n143) );
  CND2XL U1346 ( .A(n1805), .B(n835), .Z(n836) );
  CND2X1 U1347 ( .A(n834), .B(n1051), .Z(n837) );
  CND2X1 U1348 ( .A(n836), .B(n837), .Z(n1809) );
  CIVXL U1349 ( .A(n1051), .Z(n835) );
  CND2X1 U1350 ( .A(n1040), .B(n1041), .Z(n1039) );
  CND2X2 U1351 ( .A(n1093), .B(n1165), .Z(n1410) );
  CND3XL U1352 ( .A(n1086), .B(n1413), .C(n549), .Z(n1385) );
  CND3XL U1353 ( .A(n885), .B(n1413), .C(n839), .Z(n884) );
  CIVXL U1354 ( .A(n877), .Z(n885) );
  CND4XL U1355 ( .A(n884), .B(n881), .C(n883), .D(n882), .Z(n152) );
  CND3XL U1356 ( .A(n1687), .B(n1413), .C(n840), .Z(n1688) );
  CIVXL U1357 ( .A(n1684), .Z(n1687) );
  CIVXL U1358 ( .A(n1685), .Z(n1686) );
  CND4XL U1359 ( .A(n1688), .B(n1691), .C(n1689), .D(n1690), .Z(n137) );
  CNR2X1 U1360 ( .A(n1717), .B(n1192), .Z(n1144) );
  CENX1 U1361 ( .A(n1886), .B(n548), .Z(n1888) );
  CND2XL U1362 ( .A(n1891), .B(n682), .Z(n1874) );
  CND2X1 U1363 ( .A(n852), .B(n851), .Z(n845) );
  CIVXL U1364 ( .A(n845), .Z(n1169) );
  CND3XL U1365 ( .A(n846), .B(n1101), .C(n854), .Z(n853) );
  CND4XL U1366 ( .A(n846), .B(n1101), .C(n1672), .D(n1677), .Z(n1673) );
  CND2XL U1367 ( .A(n846), .B(n1164), .Z(n1163) );
  CND2XL U1368 ( .A(n846), .B(n1716), .Z(n1717) );
  CND2XL U1369 ( .A(n846), .B(n1729), .Z(n1730) );
  CND3XL U1370 ( .A(n846), .B(n1731), .C(n1729), .Z(n1725) );
  COND3XL U1371 ( .A(n847), .B(n1694), .C(n848), .D(n855), .Z(n138) );
  CND3XL U1372 ( .A(n860), .B(n1413), .C(n847), .Z(n848) );
  COND1X1 U1373 ( .A(n1911), .B(n988), .C(n849), .Z(n175) );
  COND1X1 U1374 ( .A(n1911), .B(n983), .C(n850), .Z(n179) );
  CND2IX1 U1375 ( .B(n1426), .A(n1646), .Z(n851) );
  CND2XL U1376 ( .A(n868), .B(n1426), .Z(n852) );
  CIVX2 U1377 ( .A(n1693), .Z(n854) );
  CAN2XL U1378 ( .A(n1695), .B(n1197), .Z(n860) );
  CND4XL U1379 ( .A(n1756), .B(n1758), .C(n1757), .D(n1759), .Z(n151) );
  CND3XL U1380 ( .A(n1308), .B(n1307), .C(n1309), .Z(n861) );
  CND3XL U1381 ( .A(n1308), .B(n1307), .C(n1309), .Z(n1523) );
  CMXI2X1 U1382 ( .A0(n1446), .A1(n864), .S(n546), .Z(n865) );
  CMXI2X1 U1383 ( .A0(n1444), .A1(n864), .S(n547), .Z(n1507) );
  CMXI2XL U1384 ( .A0(n1517), .A1(n865), .S(n544), .Z(n866) );
  COAN1XL U1385 ( .A(n1351), .B(n865), .C(n1193), .Z(n1349) );
  COR2X1 U1386 ( .A(n1633), .B(n866), .Z(n867) );
  CANR1XL U1387 ( .A(n1427), .B(n866), .C(n1429), .Z(n1267) );
  CND2X1 U1388 ( .A(n868), .B(n1412), .Z(n869) );
  CND2X2 U1389 ( .A(n1852), .B(n869), .Z(n878) );
  CAN2XL U1390 ( .A(n1852), .B(n869), .Z(n903) );
  CNR2X2 U1391 ( .A(n870), .B(n872), .Z(n871) );
  CNR2X1 U1392 ( .A(n927), .B(n872), .Z(n1093) );
  CND2X2 U1393 ( .A(n879), .B(n878), .Z(n873) );
  CIVX2 U1394 ( .A(n873), .Z(n880) );
  CNR2X1 U1395 ( .A(n927), .B(n873), .Z(n1407) );
  CIVX2 U1396 ( .A(n874), .Z(n1165) );
  CND2X2 U1397 ( .A(n1123), .B(n1146), .Z(n875) );
  CIVX2 U1398 ( .A(n875), .Z(n876) );
  CIVX2 U1399 ( .A(n875), .Z(n1028) );
  CND2X1 U1400 ( .A(n1098), .B(n876), .Z(n1805) );
  CAN3XL U1401 ( .A(n876), .B(n1796), .C(n1752), .Z(n1409) );
  CND3XL U1402 ( .A(n876), .B(n1796), .C(n1770), .Z(n1772) );
  CND2XL U1403 ( .A(n404), .B(n1760), .Z(n881) );
  CND2X2 U1404 ( .A(n1853), .B(n1854), .Z(n879) );
  CAOR2XL U1405 ( .A(acc[44]), .B(n1416), .C(n1195), .D(acc_a[44]), .Z(n886)
         );
  CANR1XL U1406 ( .A(n1196), .B(\C1/DATA1_44 ), .C(n886), .Z(n882) );
  CNR2X2 U1407 ( .A(n1913), .B(n887), .Z(n1891) );
  CNR2X1 U1408 ( .A(n887), .B(n893), .Z(n894) );
  CND2X1 U1409 ( .A(n888), .B(n554), .Z(n185) );
  CIVXL U1410 ( .A(n1187), .Z(n893) );
  CND2IXL U1411 ( .B(n1913), .A(n894), .Z(n891) );
  CENXL U1412 ( .A(n891), .B(n1085), .Z(n890) );
  COND4CX1 U1413 ( .A(n1927), .B(n890), .C(n892), .D(n1417), .Z(n888) );
  COND1X1 U1414 ( .A(n1911), .B(n900), .C(n895), .Z(n174) );
  COND1X1 U1415 ( .A(n1911), .B(n905), .C(n896), .Z(n178) );
  COND1XL U1416 ( .A(n898), .B(n899), .C(n547), .Z(n897) );
  CENXL U1417 ( .A(n903), .B(n904), .Z(n900) );
  CAN2XL U1418 ( .A(n1861), .B(n1860), .Z(n908) );
  CENXL U1419 ( .A(n908), .B(n909), .Z(n905) );
  CMXI2X1 U1420 ( .A0(n1790), .A1(n1078), .S(n1426), .Z(n1795) );
  CMXI2X1 U1421 ( .A0(n1467), .A1(n1466), .S(n1419), .Z(n948) );
  COR2X1 U1422 ( .A(n1633), .B(n1624), .Z(n1636) );
  CMXI2XL U1423 ( .A0(n1511), .A1(n960), .S(n1207), .Z(n911) );
  CMXI2XL U1424 ( .A0(n1481), .A1(n1551), .S(n1207), .Z(n1118) );
  CMXI2XL U1425 ( .A0(n1494), .A1(n1480), .S(n1420), .Z(n1551) );
  CMXI2X1 U1426 ( .A0(acc[23]), .A1(acc[24]), .S(n435), .Z(n1452) );
  CMXI2XL U1427 ( .A0(acc[55]), .A1(acc[54]), .S(n921), .Z(n1441) );
  CND2IX1 U1428 ( .B(n540), .A(n1567), .Z(n1315) );
  CMXI2X1 U1429 ( .A0(n1652), .A1(n1639), .S(n1423), .Z(n1789) );
  CND4X1 U1430 ( .A(n1155), .B(n1152), .C(n1154), .D(n1153), .Z(n139) );
  CMXI2X1 U1431 ( .A0(n1506), .A1(n1507), .S(n1207), .Z(n1562) );
  CIVDX2 U1432 ( .A(n544), .Z0(n1203), .Z1(n1204) );
  CAN2X1 U1433 ( .A(n1860), .B(n1861), .Z(n1048) );
  COR2XL U1434 ( .A(n1633), .B(n1562), .Z(n920) );
  CNR2XL U1435 ( .A(n1673), .B(n1192), .Z(n1676) );
  CND3XL U1436 ( .A(n961), .B(n1349), .C(n1350), .Z(n972) );
  CMXI2X1 U1437 ( .A0(n1563), .A1(n1562), .S(ho_2[5]), .Z(n1564) );
  CMXI2XL U1438 ( .A0(n1578), .A1(n1577), .S(n1424), .Z(n1580) );
  CIVX8 U1439 ( .A(n921), .Z(n922) );
  CMXI2X1 U1440 ( .A0(n1453), .A1(n1452), .S(n1419), .Z(n1555) );
  CIVX8 U1441 ( .A(n546), .Z(n1420) );
  CANR1X1 U1442 ( .A(\DP_OP_14_298_9081/n95 ), .B(\DP_OP_14_298_9081/n2 ), .C(
        \DP_OP_14_298_9081/n96 ), .Z(\DP_OP_14_298_9081/n94 ) );
  COAN1XL U1443 ( .A(n1310), .B(n1507), .C(n1193), .Z(n1307) );
  CMXI2X1 U1444 ( .A0(n1105), .A1(n1487), .S(n923), .Z(n1106) );
  CMXI2XL U1445 ( .A0(n1575), .A1(n1550), .S(n1419), .Z(n1556) );
  CND2IXL U1446 ( .B(n686), .A(n1277), .Z(n1276) );
  CMXI2X1 U1447 ( .A0(n1112), .A1(n1504), .S(n1204), .Z(n1612) );
  CMXI2XL U1448 ( .A0(acc[13]), .A1(n1095), .S(n922), .Z(n1554) );
  CND2IXL U1449 ( .B(n923), .A(n963), .Z(n980) );
  CNR2XL U1450 ( .A(n680), .B(acc_a[38]), .Z(\DP_OP_14_298_9081/n252 ) );
  CMX2XL U1451 ( .A0(n415), .A1(n465), .S(ho_2[2]), .Z(n928) );
  CIVXL U1452 ( .A(n928), .Z(n929) );
  CMXI2X1 U1453 ( .A0(n1640), .A1(n1639), .S(ho_2[2]), .Z(n1723) );
  CND2IX1 U1454 ( .B(n686), .A(n1229), .Z(n1230) );
  CANR1X1 U1455 ( .A(n1421), .B(n1596), .C(n1412), .Z(n976) );
  CNR2IX2 U1456 ( .B(n1407), .A(n1858), .Z(n1851) );
  CND3X2 U1457 ( .A(n1289), .B(n1290), .C(n1291), .Z(n1515) );
  COND1XL U1458 ( .A(n923), .B(n1529), .C(n540), .Z(n935) );
  CND3XL U1459 ( .A(n1003), .B(n1002), .C(n1784), .Z(n936) );
  CND2XL U1460 ( .A(n681), .B(acc_a[38]), .Z(\DP_OP_14_298_9081/n253 ) );
  CND2IX1 U1461 ( .B(n1633), .A(n938), .Z(n946) );
  CMX2XL U1462 ( .A0(n1478), .A1(n1477), .S(n1424), .Z(n938) );
  CMXI2X1 U1463 ( .A0(n1515), .A1(n1484), .S(n1423), .Z(n1590) );
  CND2X1 U1464 ( .A(n1131), .B(n1130), .Z(n1115) );
  CNIVXL U1465 ( .A(n1106), .Z(n1078) );
  CND2IX1 U1466 ( .B(n1425), .A(n1645), .Z(n1223) );
  CMXI2X1 U1467 ( .A0(n1595), .A1(n1596), .S(n542), .Z(n1121) );
  CMXI2XL U1468 ( .A0(n1478), .A1(n1477), .S(n1424), .Z(n939) );
  CND2IXL U1469 ( .B(n1425), .A(n1077), .Z(n940) );
  CND2IXL U1470 ( .B(n1428), .A(n1603), .Z(n1254) );
  CND2XL U1471 ( .A(n1160), .B(n1159), .Z(n941) );
  CMXI2X1 U1472 ( .A0(n1482), .A1(n1483), .S(n1207), .Z(n1528) );
  COND1XL U1473 ( .A(n1911), .B(n1166), .C(n1167), .Z(n158) );
  CND2XL U1474 ( .A(n1171), .B(n1172), .Z(n1166) );
  CND3XL U1475 ( .A(n1873), .B(n1187), .C(n1875), .Z(n942) );
  CND2XL U1476 ( .A(n1891), .B(n943), .Z(n1866) );
  CIVXL U1477 ( .A(n942), .Z(n943) );
  CENXL U1478 ( .A(n1050), .B(n1363), .Z(n1360) );
  CMXI2X1 U1479 ( .A0(n1518), .A1(n1526), .S(n543), .Z(n1246) );
  CND2X2 U1480 ( .A(n1282), .B(n1283), .Z(n1922) );
  CNR2X1 U1481 ( .A(n1126), .B(n1127), .Z(n1125) );
  CMXI2XL U1482 ( .A0(n1467), .A1(n1466), .S(n1419), .Z(n947) );
  CND2XL U1483 ( .A(n1108), .B(n1107), .Z(n1574) );
  CENXL U1484 ( .A(n996), .B(n949), .Z(n993) );
  CND2IX1 U1485 ( .B(n1426), .A(n1058), .Z(n1103) );
  CND2XL U1486 ( .A(n1806), .B(n1804), .Z(n950) );
  CND2XL U1487 ( .A(n941), .B(n1804), .Z(n951) );
  CND2X1 U1488 ( .A(n1631), .B(n1423), .Z(n952) );
  CND2IX2 U1489 ( .B(n1426), .A(n677), .Z(n1336) );
  CMXI2XL U1490 ( .A0(n947), .A1(n960), .S(n545), .Z(n955) );
  CMXI2XL U1491 ( .A0(n948), .A1(n960), .S(n545), .Z(n1579) );
  CND2IXL U1492 ( .B(n1425), .A(n1538), .Z(n1260) );
  CND2IXL U1493 ( .B(n541), .A(n1538), .Z(n1324) );
  CNR2XL U1494 ( .A(n1813), .B(n1911), .Z(n1814) );
  CANR1X1 U1495 ( .A(\DP_OP_14_298_9081/n176 ), .B(\DP_OP_14_298_9081/n163 ), 
        .C(\DP_OP_14_298_9081/n164 ), .Z(\DP_OP_14_298_9081/n158 ) );
  CNR2IX2 U1496 ( .B(n1723), .A(n1726), .Z(n1706) );
  CND3XL U1497 ( .A(n1005), .B(n1007), .C(n1009), .Z(n134) );
  CND2XL U1498 ( .A(n926), .B(acc_a[62]), .Z(\DP_OP_14_298_9081/n73 ) );
  CNR2XL U1499 ( .A(n926), .B(acc_a[62]), .Z(\DP_OP_14_298_9081/n72 ) );
  CMXI2X1 U1500 ( .A0(acc[44]), .A1(n309), .S(n1418), .Z(n1449) );
  CMXI2X1 U1501 ( .A0(acc[36]), .A1(n944), .S(n922), .Z(n1444) );
  CMXI2X1 U1502 ( .A0(acc[26]), .A1(acc[27]), .S(n1418), .Z(n1443) );
  CMXI2X1 U1503 ( .A0(acc[19]), .A1(acc[20]), .S(n922), .Z(n1480) );
  CMXI2X1 U1504 ( .A0(acc[27]), .A1(acc[28]), .S(n922), .Z(n1460) );
  CMXI2X1 U1505 ( .A0(acc[29]), .A1(acc[30]), .S(n922), .Z(n1455) );
  CMXI2X1 U1506 ( .A0(n958), .A1(n1468), .S(n1420), .Z(n960) );
  CMXI2X1 U1507 ( .A0(n1469), .A1(n958), .S(n1420), .Z(n1504) );
  CMXI2XL U1508 ( .A0(n1511), .A1(n960), .S(n1207), .Z(n962) );
  CND3XL U1509 ( .A(n1349), .B(n961), .C(n1350), .Z(n1054) );
  COR2X1 U1510 ( .A(n1633), .B(n911), .Z(n1529) );
  CND2IXL U1511 ( .B(n1422), .A(n963), .Z(n1228) );
  CMXI2X1 U1512 ( .A0(n1520), .A1(n972), .S(n1422), .Z(n964) );
  CND2IXL U1513 ( .B(n1426), .A(n964), .Z(n975) );
  CND2IXL U1514 ( .B(n541), .A(n964), .Z(n1040) );
  CMXI2XL U1515 ( .A0(n1246), .A1(n964), .S(n1425), .Z(n1848) );
  CND2X1 U1516 ( .A(n980), .B(n981), .Z(n965) );
  CND2X1 U1517 ( .A(n1179), .B(n965), .Z(n966) );
  CND2XL U1518 ( .A(n940), .B(n965), .Z(n1052) );
  CND2X2 U1519 ( .A(n966), .B(n967), .Z(n968) );
  CND2XL U1520 ( .A(n1881), .B(n966), .Z(n1231) );
  CND2X1 U1521 ( .A(n975), .B(n974), .Z(n967) );
  CIVXL U1522 ( .A(n967), .Z(n1373) );
  CNR2X2 U1523 ( .A(n1237), .B(n968), .Z(n1187) );
  CND3XL U1524 ( .A(n1891), .B(n1085), .C(n1187), .Z(n1343) );
  CIVX2 U1525 ( .A(n969), .Z(n1335) );
  CAN2XL U1526 ( .A(n1012), .B(n1010), .Z(n970) );
  CND3XL U1527 ( .A(n1011), .B(n970), .C(n1013), .Z(n141) );
  CND2IX1 U1528 ( .B(n1423), .A(n1619), .Z(n971) );
  COND2XL U1529 ( .A(n540), .B(n1655), .C(n1218), .D(n1219), .Z(n973) );
  COR2X1 U1530 ( .A(n1773), .B(n973), .Z(n1122) );
  CND2IX1 U1531 ( .B(n1421), .A(n1586), .Z(n977) );
  CANR1X1 U1532 ( .A(n1422), .B(n1594), .C(n541), .Z(n978) );
  CANR1XL U1533 ( .A(n1276), .B(n1275), .C(n1422), .Z(n979) );
  CND2IX1 U1534 ( .B(n979), .A(n978), .Z(n1132) );
  CANR1X1 U1535 ( .A(n923), .B(n1588), .C(n1411), .Z(n981) );
  CND2XL U1536 ( .A(n1098), .B(n1863), .Z(n987) );
  CENXL U1537 ( .A(n986), .B(n987), .Z(n983) );
  CND2XL U1538 ( .A(n1098), .B(n1856), .Z(n992) );
  CENXL U1539 ( .A(n991), .B(n992), .Z(n988) );
  CNR3XL U1540 ( .A(n1791), .B(n1785), .C(n1787), .Z(n997) );
  CAOR2XL U1541 ( .A(acc[40]), .B(n1416), .C(n1195), .D(acc_a[40]), .Z(n995)
         );
  CND3XL U1542 ( .A(n969), .B(n912), .C(n997), .Z(n996) );
  CANR1XL U1543 ( .A(n1196), .B(\C1/DATA1_40 ), .C(n995), .Z(n994) );
  COND1X1 U1544 ( .A(n1911), .B(n993), .C(n994), .Z(n156) );
  CND2IX1 U1545 ( .B(n1001), .A(n541), .Z(n1325) );
  CND2XL U1546 ( .A(n1001), .B(n1426), .Z(n1003) );
  CNR2XL U1547 ( .A(n1122), .B(n936), .Z(n1057) );
  CMXI2XL U1548 ( .A0(n1450), .A1(n1446), .S(n546), .Z(n998) );
  CMXI2XL U1549 ( .A0(n1490), .A1(n998), .S(n1204), .Z(n1104) );
  COR2X1 U1550 ( .A(n1633), .B(n1104), .Z(n1105) );
  CND2X1 U1551 ( .A(n1521), .B(n1422), .Z(n1000) );
  CND2X1 U1552 ( .A(n1105), .B(n1423), .Z(n999) );
  CND2X1 U1553 ( .A(n999), .B(n1000), .Z(n1001) );
  CAOR2XL U1554 ( .A(n926), .B(n1416), .C(n1195), .D(acc_a[62]), .Z(n1008) );
  CANR1XL U1555 ( .A(n1196), .B(\C1/DATA1_62 ), .C(n1008), .Z(n1004) );
  CND4XL U1556 ( .A(n1247), .B(n1413), .C(n1197), .D(n1671), .Z(n1007) );
  CAOR2XL U1557 ( .A(acc[55]), .B(n1416), .C(n1195), .D(acc_a[55]), .Z(n1014)
         );
  CANR1XL U1558 ( .A(n1196), .B(\C1/DATA1_55 ), .C(n1014), .Z(n1010) );
  CND4XL U1559 ( .A(n1248), .B(n1413), .C(n1197), .D(n1704), .Z(n1013) );
  CND2IXL U1560 ( .B(n1426), .A(n1106), .Z(n1015) );
  CND2X1 U1561 ( .A(n1015), .B(n1016), .Z(n1182) );
  CMXI2X1 U1562 ( .A0(n1521), .A1(n1631), .S(n1422), .Z(n1017) );
  CMXI2XL U1563 ( .A0(n1743), .A1(n1017), .S(n1426), .Z(n1761) );
  CND2X2 U1564 ( .A(n1019), .B(n1020), .Z(n1111) );
  CND2IX1 U1565 ( .B(n1021), .A(n1110), .Z(n1019) );
  CND2IX2 U1566 ( .B(n543), .A(n1641), .Z(n1020) );
  CNR2XL U1567 ( .A(n1552), .B(n1633), .Z(n1024) );
  CND2XL U1568 ( .A(n1024), .B(n685), .Z(n1023) );
  COND1X1 U1569 ( .A(n685), .B(n1529), .C(n1023), .Z(n1025) );
  CND2IX1 U1570 ( .B(n1426), .A(n1025), .Z(n1042) );
  CND2X2 U1571 ( .A(n1039), .B(n1038), .Z(n1026) );
  CIVX2 U1572 ( .A(n1027), .Z(n1123) );
  CIVX2 U1573 ( .A(n1028), .Z(n1191) );
  CMXI2X1 U1574 ( .A0(n1471), .A1(n1472), .S(n546), .Z(n1483) );
  CMXI2X1 U1575 ( .A0(n1483), .A1(n1477), .S(n544), .Z(n1552) );
  COAN1X1 U1576 ( .A(n1204), .B(n1556), .C(n1035), .Z(n1033) );
  CND2IX1 U1577 ( .B(n1203), .A(n1036), .Z(n1032) );
  CAOR1X1 U1578 ( .A(n1419), .B(n1583), .C(n1037), .Z(n1036) );
  COR2XL U1579 ( .A(n1031), .B(n1229), .Z(n1030) );
  CND2IX1 U1580 ( .B(n1425), .A(n1246), .Z(n1041) );
  CND2IXL U1581 ( .B(n541), .A(n1846), .Z(n1043) );
  CND2X1 U1582 ( .A(n1043), .B(n1042), .Z(n1038) );
  CNR2X2 U1583 ( .A(n1813), .B(n1820), .Z(n1044) );
  CNR2IXL U1584 ( .B(n1128), .A(n1555), .Z(n1127) );
  CAN2XL U1585 ( .A(n1894), .B(n1895), .Z(n1908) );
  CMXI2X1 U1586 ( .A0(n1524), .A1(n1499), .S(n1280), .Z(n1500) );
  CMXI2XL U1587 ( .A0(n1452), .A1(n1461), .S(n1419), .Z(n1495) );
  CMXI2XL U1588 ( .A0(n1505), .A1(n1509), .S(n545), .Z(n1046) );
  CMXI2XL U1589 ( .A0(n1505), .A1(n1509), .S(n545), .Z(n1630) );
  CND2IXL U1590 ( .B(n1280), .A(n1630), .Z(n1241) );
  CND2IXL U1591 ( .B(n1421), .A(n1591), .Z(n1262) );
  CNR2XL U1592 ( .A(n1913), .B(n1906), .Z(n1907) );
  CNR2X1 U1593 ( .A(n1048), .B(n986), .Z(n1406) );
  CND2X2 U1594 ( .A(n1863), .B(n1406), .Z(n1858) );
  CMXI2XL U1595 ( .A0(n1572), .A1(n1571), .S(n1419), .Z(n1274) );
  CMXI2XL U1596 ( .A0(n1571), .A1(n1569), .S(n1419), .Z(n1561) );
  CND2X2 U1597 ( .A(n1408), .B(n409), .Z(n1913) );
  CMXI2XL U1598 ( .A0(n1583), .A1(n1582), .S(n1419), .Z(n1288) );
  CIVXL U1599 ( .A(n1803), .Z(n1049) );
  CMXI2X1 U1600 ( .A0(n1461), .A1(n1460), .S(n1420), .Z(n1481) );
  CND2IXL U1601 ( .B(n543), .A(n1529), .Z(n1221) );
  CIVXL U1602 ( .A(n1804), .Z(n1050) );
  CNIVX1 U1603 ( .A(n941), .Z(n1051) );
  CND2IX1 U1604 ( .B(n1194), .A(n1500), .Z(n1594) );
  CNR2X1 U1605 ( .A(n1730), .B(n307), .Z(n1158) );
  CND2X1 U1606 ( .A(n1263), .B(n1264), .Z(n1585) );
  COR2X1 U1607 ( .A(n1633), .B(n1626), .Z(n1637) );
  CND2IX1 U1608 ( .B(n1203), .A(n1482), .Z(n1604) );
  CMXI2XL U1609 ( .A0(n465), .A1(n1652), .S(n543), .Z(n1053) );
  CMXI2XL U1610 ( .A0(acc[1]), .A1(acc[2]), .S(n922), .Z(n1583) );
  CMXI2XL U1611 ( .A0(acc[6]), .A1(acc[7]), .S(n922), .Z(n1569) );
  CMXI2XL U1612 ( .A0(acc[4]), .A1(acc[5]), .S(n922), .Z(n1571) );
  CMXI2XL U1613 ( .A0(acc[8]), .A1(acc[9]), .S(n922), .Z(n1568) );
  CNR2X2 U1614 ( .A(n922), .B(n1435), .Z(n1456) );
  CANR1X1 U1615 ( .A(n1421), .B(n1593), .C(n1411), .Z(n1261) );
  CAN2XL U1616 ( .A(n1863), .B(n1406), .Z(n1056) );
  CND2X2 U1617 ( .A(n1328), .B(n1329), .Z(n1794) );
  CDLY1XL U1618 ( .A(n1773), .Z(n1072) );
  CMXI2X1 U1619 ( .A0(n1479), .A1(n946), .S(n685), .Z(n1058) );
  COND2XL U1620 ( .A(n540), .B(n1655), .C(n935), .D(n1218), .Z(n1059) );
  CND2IXL U1621 ( .B(n542), .A(n1491), .Z(n1352) );
  CND3XL U1622 ( .A(n1156), .B(n1413), .C(n1060), .Z(n1155) );
  CMXI2X1 U1623 ( .A0(n1508), .A1(n1534), .S(n544), .Z(n1243) );
  CNR2XL U1624 ( .A(n1720), .B(n1722), .Z(n1716) );
  CMXI2X1 U1625 ( .A0(n1491), .A1(n1510), .S(ho_2[2]), .Z(n1857) );
  CMXI2XL U1626 ( .A0(n1506), .A1(n1505), .S(n1206), .Z(n1535) );
  CND2IX1 U1627 ( .B(n1611), .A(n1035), .Z(n1110) );
  CANR1X1 U1628 ( .A(n686), .B(n1611), .C(n1194), .Z(n1263) );
  CND2X2 U1629 ( .A(n1226), .B(n1225), .Z(n1875) );
  CND2X1 U1630 ( .A(n1227), .B(n1228), .Z(n1225) );
  CND2XL U1631 ( .A(n1874), .B(n1066), .Z(n1067) );
  CND2XL U1632 ( .A(n1065), .B(n1875), .Z(n1068) );
  CND2X1 U1633 ( .A(n1067), .B(n1068), .Z(n1879) );
  CIVXL U1634 ( .A(n1874), .Z(n1065) );
  CIVXL U1635 ( .A(n1875), .Z(n1066) );
  CND4X1 U1636 ( .A(n1775), .B(n1777), .C(n1776), .D(n1778), .Z(n154) );
  CIVXL U1637 ( .A(n1708), .Z(n1711) );
  CMXI2XL U1638 ( .A0(n1569), .A1(n1568), .S(n1419), .Z(n1269) );
  CMXI2XL U1639 ( .A0(n1565), .A1(n1531), .S(n545), .Z(n1532) );
  CMXI2XL U1640 ( .A0(n1321), .A1(n1565), .S(n1203), .Z(n1320) );
  CND2X1 U1641 ( .A(n1479), .B(n685), .Z(n1073) );
  CND2X2 U1642 ( .A(n1512), .B(n543), .Z(n1074) );
  CND2X2 U1643 ( .A(n1073), .B(n1074), .Z(n1075) );
  CND2IX1 U1644 ( .B(n1411), .A(n1628), .Z(n1328) );
  CND2X2 U1645 ( .A(n1628), .B(n1411), .Z(n1853) );
  CMXI2XL U1646 ( .A0(n1515), .A1(n1527), .S(n1422), .Z(n1077) );
  CMXI2X1 U1647 ( .A0(n1462), .A1(n1463), .S(n546), .Z(n1478) );
  CAN2XL U1648 ( .A(n1646), .B(n1425), .Z(n1708) );
  CMX2XL U1649 ( .A0(n1660), .A1(n666), .S(n1426), .Z(n1081) );
  CND2X1 U1650 ( .A(n1567), .B(n1426), .Z(n1084) );
  CND2X2 U1651 ( .A(n1696), .B(n1656), .Z(n1693) );
  CNR2X2 U1652 ( .A(n1704), .B(n1701), .Z(n1696) );
  CND4XL U1653 ( .A(n1409), .B(n1197), .C(n1252), .D(n1413), .Z(n1756) );
  CMXI2XL U1654 ( .A0(n1269), .A1(n1570), .S(n1206), .Z(n1268) );
  CNR3X1 U1655 ( .A(n1913), .B(n1906), .C(n1908), .Z(n1901) );
  CEOXL U1656 ( .A(n1908), .B(n1907), .Z(n1912) );
  CND2IXL U1657 ( .B(n1913), .A(n1080), .Z(n1882) );
  CANR1X1 U1658 ( .A(n1280), .B(n1281), .C(n1429), .Z(n1278) );
  CENXL U1659 ( .A(n1314), .B(n1079), .Z(n1311) );
  CND2XL U1660 ( .A(n1261), .B(n1262), .Z(n1259) );
  COND1X1 U1661 ( .A(n1422), .B(n1518), .C(n540), .Z(n1245) );
  CND2X2 U1662 ( .A(n1149), .B(n1148), .Z(n1236) );
  CND2IX1 U1663 ( .B(n540), .A(n1061), .Z(n1148) );
  CAN2XL U1664 ( .A(n1657), .B(n1425), .Z(n1692) );
  COND1X1 U1665 ( .A(n1423), .B(n1529), .C(n540), .Z(n1219) );
  CMXI2X1 U1666 ( .A0(n1641), .A1(n1642), .S(n542), .Z(n1082) );
  CMXI2X1 U1667 ( .A0(n1641), .A1(n1642), .S(n542), .Z(n1643) );
  CND2IXL U1668 ( .B(n1280), .A(n1605), .Z(n1302) );
  CMXI2XL U1669 ( .A0(n1530), .A1(n1495), .S(n1206), .Z(n1499) );
  CIVX2 U1670 ( .A(n1079), .Z(n1864) );
  CND2X2 U1671 ( .A(n1249), .B(n1250), .Z(n1629) );
  CAN2X1 U1672 ( .A(n1865), .B(n1864), .Z(n1863) );
  CNR2XL U1673 ( .A(n1380), .B(n307), .Z(n1086) );
  CNR2X2 U1674 ( .A(n1334), .B(n1917), .Z(n1408) );
  CMXI2XL U1675 ( .A0(n1322), .A1(n1572), .S(n1419), .Z(n1321) );
  CANR1X1 U1676 ( .A(n1422), .B(n1598), .C(n1411), .Z(n1227) );
  CIVXL U1677 ( .A(n1906), .Z(n1088) );
  CIVX2 U1678 ( .A(n1335), .Z(n1414) );
  CND2IXL U1679 ( .B(n1616), .A(n1650), .Z(n1617) );
  CNR2X2 U1680 ( .A(n1722), .B(n1719), .Z(n1707) );
  CND2X1 U1681 ( .A(n1232), .B(n1233), .Z(n1595) );
  CND2XL U1682 ( .A(n1090), .B(n1867), .Z(n1091) );
  CND2XL U1683 ( .A(n1866), .B(n1089), .Z(n1092) );
  CND2XL U1684 ( .A(n1091), .B(n1092), .Z(n1871) );
  CIVXL U1685 ( .A(n1867), .Z(n1089) );
  CIVXL U1686 ( .A(n1866), .Z(n1090) );
  COND4CXL U1687 ( .A(n1872), .B(n1871), .C(n1870), .D(n1869), .Z(n182) );
  CND2X2 U1688 ( .A(n1867), .B(n1875), .Z(n1145) );
  CND2X2 U1689 ( .A(n1326), .B(n1327), .Z(n1820) );
  CIVXL U1690 ( .A(n1222), .Z(n1399) );
  CND2XL U1691 ( .A(n302), .B(n1741), .Z(n1097) );
  CND2IXL U1692 ( .B(n1508), .A(n1293), .Z(n1309) );
  CMXI2XL U1693 ( .A0(n1560), .A1(n1534), .S(n545), .Z(n1536) );
  CMXI2XL U1694 ( .A0(n1561), .A1(n1560), .S(n1203), .Z(n1563) );
  CND2IXL U1695 ( .B(n1747), .A(n1748), .Z(n1296) );
  CMXI2XL U1696 ( .A0(n1446), .A1(n1450), .S(n547), .Z(n1099) );
  CND2XL U1697 ( .A(n1853), .B(n1854), .Z(n1855) );
  CAN2XL U1698 ( .A(n933), .B(n1197), .Z(n1390) );
  CNR2XL U1699 ( .A(n933), .B(n1911), .Z(n1394) );
  COR2X1 U1700 ( .A(n1633), .B(n1528), .Z(n1638) );
  CIVX2 U1701 ( .A(n1702), .Z(n1100) );
  CIVX2 U1702 ( .A(n1100), .Z(n1101) );
  CNR2XL U1703 ( .A(n1072), .B(n1911), .Z(n1771) );
  CMXI2X1 U1704 ( .A0(acc[59]), .A1(acc[60]), .S(n922), .Z(n1464) );
  CND2XL U1705 ( .A(n1102), .B(n1426), .Z(n1224) );
  CND2X1 U1706 ( .A(n1103), .B(n1116), .Z(n1862) );
  CMXI2X1 U1707 ( .A0(n1470), .A1(n1469), .S(n1420), .Z(n1477) );
  CND2IX1 U1708 ( .B(n543), .A(n1595), .Z(n1108) );
  CMXI2X1 U1709 ( .A0(n1480), .A1(n1453), .S(n1420), .Z(n1109) );
  CMXI2XL U1710 ( .A0(n1558), .A1(n1109), .S(n545), .Z(n1277) );
  CIVX2 U1711 ( .A(n1111), .Z(n1788) );
  CMXI2X1 U1712 ( .A0(n1466), .A1(n1470), .S(n1419), .Z(n1492) );
  CMXI2X1 U1713 ( .A0(n1492), .A1(n1498), .S(n1424), .Z(n1611) );
  CMXI2X1 U1714 ( .A0(n1471), .A1(n1459), .S(n547), .Z(n1112) );
  CND2IX1 U1715 ( .B(n1426), .A(n1082), .Z(n1114) );
  CND2IX1 U1716 ( .B(n1411), .A(n1501), .Z(n1113) );
  CND2X2 U1717 ( .A(n1115), .B(n541), .Z(n1282) );
  CND3X2 U1718 ( .A(n1131), .B(n1130), .C(n1426), .Z(n1116) );
  CND2IX1 U1719 ( .B(n1194), .A(n1117), .Z(n1598) );
  CND2IX1 U1720 ( .B(n1426), .A(n1597), .Z(n1120) );
  CND2X1 U1721 ( .A(n1119), .B(n1120), .Z(n1867) );
  CND2XL U1722 ( .A(n1426), .B(n1121), .Z(n1119) );
  CND3XL U1723 ( .A(n1851), .B(n1076), .C(n1832), .Z(n1836) );
  CAN3XL U1724 ( .A(n1076), .B(n945), .C(n1810), .Z(n1201) );
  CAN2XL U1725 ( .A(n1076), .B(n945), .Z(n1202) );
  CND2IX1 U1726 ( .B(n686), .A(n545), .Z(n1129) );
  CND2IXL U1727 ( .B(n1280), .A(n1626), .Z(n1124) );
  CND2X1 U1728 ( .A(n1124), .B(n1125), .Z(n1484) );
  CND2IX1 U1729 ( .B(n1423), .A(n1484), .Z(n1130) );
  CND2IX1 U1730 ( .B(n1426), .A(n1134), .Z(n1133) );
  COR2X1 U1731 ( .A(n1633), .B(n1579), .Z(n1479) );
  CIVXL U1732 ( .A(n927), .Z(n1185) );
  CND3X1 U1733 ( .A(n1141), .B(n1140), .C(n1135), .Z(n144) );
  CND2IX1 U1734 ( .B(n1422), .A(n1589), .Z(n1138) );
  CND2IXL U1735 ( .B(n540), .A(n934), .Z(n1137) );
  CND2X1 U1736 ( .A(n1137), .B(n1136), .Z(n1902) );
  CND2X1 U1737 ( .A(n1138), .B(n1139), .Z(n1136) );
  CAOR2XL U1738 ( .A(acc[52]), .B(n1416), .C(n1195), .D(acc_a[52]), .Z(n1143)
         );
  CIVXL U1739 ( .A(n1144), .Z(n1142) );
  CND4XL U1740 ( .A(n1144), .B(n1413), .C(n1197), .D(n1719), .Z(n1141) );
  CND2X1 U1741 ( .A(n1142), .B(n1718), .Z(n1140) );
  CND2IXL U1742 ( .B(n1421), .A(n1585), .Z(n1151) );
  CND3X1 U1743 ( .A(n1150), .B(n1151), .C(n540), .Z(n1149) );
  CAOR2XL U1744 ( .A(n841), .B(n1416), .C(n1195), .D(acc_a[57]), .Z(n1157) );
  CIVXL U1745 ( .A(n1698), .Z(n1156) );
  CND2XL U1746 ( .A(n1698), .B(n1697), .Z(n1152) );
  CANR1XL U1747 ( .A(n1196), .B(\C1/DATA1_57 ), .C(n1157), .Z(n1153) );
  CND2X2 U1748 ( .A(n1160), .B(n1159), .Z(n1806) );
  CND2IX1 U1749 ( .B(n1426), .A(n1723), .Z(n1160) );
  CND2IX1 U1750 ( .B(n541), .A(n1643), .Z(n1159) );
  CND2X2 U1751 ( .A(n1806), .B(n1804), .Z(n1162) );
  CIVX2 U1752 ( .A(n1162), .Z(n1161) );
  CAN2XL U1753 ( .A(n1702), .B(n1677), .Z(n1164) );
  CNR2X1 U1754 ( .A(n1163), .B(n307), .Z(n1680) );
  CIVXL U1755 ( .A(n1792), .Z(n1170) );
  CAOR2XL U1756 ( .A(n681), .B(n1416), .C(n1195), .D(acc_a[38]), .Z(n1168) );
  CND2XL U1757 ( .A(n406), .B(n1169), .Z(n1172) );
  CND2XL U1758 ( .A(n1170), .B(n1047), .Z(n1171) );
  CANR1XL U1759 ( .A(n1196), .B(\C1/DATA1_38 ), .C(n1168), .Z(n1167) );
  CND2XL U1760 ( .A(n1098), .B(n1183), .Z(n1178) );
  CENXL U1761 ( .A(n1178), .B(n1177), .Z(n1173) );
  COND1X1 U1762 ( .A(n1911), .B(n1173), .C(n1174), .Z(n173) );
  CND2IXL U1763 ( .B(n1425), .A(n1846), .Z(n1179) );
  CND3X1 U1764 ( .A(n1677), .B(n1702), .C(n1180), .Z(n1669) );
  CNR2X1 U1765 ( .A(n1181), .B(n1191), .Z(n1247) );
  CIVX4 U1766 ( .A(ho_2[5]), .Z(n1428) );
  CENXL U1767 ( .A(n1897), .B(n1896), .Z(n1900) );
  COND3XL U1768 ( .A(n1395), .B(n1387), .C(n1388), .D(n1389), .Z(n162) );
  CND2XL U1769 ( .A(n1395), .B(n1390), .Z(n1388) );
  CENXL U1770 ( .A(n1342), .B(n1343), .Z(n1338) );
  COND3XL U1771 ( .A(n1395), .B(n1205), .C(n1354), .D(n1355), .Z(n160) );
  CND2XL U1772 ( .A(n1395), .B(n1356), .Z(n1354) );
  CND4XL U1773 ( .A(n1819), .B(n1817), .C(n1818), .D(n1816), .Z(n166) );
  CND2X2 U1774 ( .A(n1270), .B(n1425), .Z(n1239) );
  CMXI2XL U1775 ( .A0(n1274), .A1(n1573), .S(n1203), .Z(n1273) );
  CMXI2XL U1776 ( .A0(n1573), .A1(n1541), .S(n545), .Z(n1543) );
  COND1X1 U1777 ( .A(n1911), .B(n1801), .C(n1800), .Z(n161) );
  CND2XL U1778 ( .A(n1267), .B(n1266), .Z(n1587) );
  CMX2XL U1779 ( .A0(n1082), .A1(n1501), .S(n1425), .Z(n1865) );
  CND2XL U1780 ( .A(n1415), .B(n1771), .Z(n1776) );
  COND1X1 U1781 ( .A(n1911), .B(n1740), .C(n1739), .Z(n149) );
  COND1X1 U1782 ( .A(n1911), .B(n1783), .C(n1782), .Z(n155) );
  CND2XL U1783 ( .A(n1772), .B(n1771), .Z(n1777) );
  CNR2X1 U1784 ( .A(n1858), .B(n1186), .Z(n1856) );
  CMXI2X1 U1785 ( .A0(n1497), .A1(n1498), .S(n1207), .Z(n1524) );
  CNR2IX2 U1786 ( .B(n1407), .A(n1858), .Z(n1183) );
  COND1X1 U1787 ( .A(n1911), .B(n1845), .C(n1844), .Z(n169) );
  COND1X1 U1788 ( .A(n1911), .B(n1768), .C(n1767), .Z(n153) );
  COND1X1 U1789 ( .A(n1911), .B(n1311), .C(n1312), .Z(n180) );
  COND3XL U1790 ( .A(n1413), .B(n1829), .C(n1828), .D(n1827), .Z(n167) );
  CND4XL U1791 ( .A(n1821), .B(n1414), .C(n1197), .D(n1820), .Z(n1828) );
  CIVX2 U1792 ( .A(n1335), .Z(n1413) );
  COND1X1 U1793 ( .A(n1911), .B(n1360), .C(n1361), .Z(n164) );
  CND2IXL U1794 ( .B(n1683), .A(n1415), .Z(n1689) );
  CND2XL U1795 ( .A(n876), .B(n1746), .Z(n1748) );
  COND3XL U1796 ( .A(n1748), .B(n1295), .C(n1296), .D(n1297), .Z(n150) );
  CND2XL U1797 ( .A(n1413), .B(n1300), .Z(n1295) );
  CMXI2XL U1798 ( .A0(acc[2]), .A1(acc[3]), .S(n922), .Z(n1572) );
  COND3XL U1799 ( .A(n1413), .B(n1840), .C(n1839), .D(n1838), .Z(n168) );
  CND4XL U1800 ( .A(n1834), .B(n1414), .C(n1197), .D(n1833), .Z(n1839) );
  CIVXL U1801 ( .A(n1185), .Z(n1186) );
  CNR2XL U1802 ( .A(n1725), .B(n306), .Z(n1727) );
  CND2IXL U1803 ( .B(n1683), .A(n1684), .Z(n1691) );
  COND1X1 U1804 ( .A(n1911), .B(n1396), .C(n1397), .Z(n172) );
  COR2X1 U1805 ( .A(n1045), .B(acc_a[61]), .Z(n1190) );
  CIVX2 U1806 ( .A(\DP_OP_14_298_9081/n427 ), .Z(\DP_OP_14_298_9081/n426 ) );
  CIVXL U1807 ( .A(\DP_OP_14_298_9081/n2 ), .Z(\DP_OP_14_298_9081/n290 ) );
  CIVXL U1808 ( .A(\DP_OP_14_298_9081/n342 ), .Z(\DP_OP_14_298_9081/n340 ) );
  CIVXL U1809 ( .A(\DP_OP_14_298_9081/n321 ), .Z(\DP_OP_14_298_9081/n319 ) );
  CIVXL U1810 ( .A(\DP_OP_14_298_9081/n3 ), .Z(\DP_OP_14_298_9081/n184 ) );
  CIVXL U1811 ( .A(\DP_OP_14_298_9081/n240 ), .Z(\DP_OP_14_298_9081/n242 ) );
  CIVXL U1812 ( .A(\DP_OP_14_298_9081/n1 ), .Z(\DP_OP_14_298_9081/n381 ) );
  CIVXL U1813 ( .A(\DP_OP_14_298_9081/n218 ), .Z(\DP_OP_14_298_9081/n216 ) );
  CIVXL U1814 ( .A(\DP_OP_14_298_9081/n214 ), .Z(\DP_OP_14_298_9081/n212 ) );
  CIVXL U1815 ( .A(\DP_OP_14_298_9081/n361 ), .Z(\DP_OP_14_298_9081/n360 ) );
  CIVXL U1816 ( .A(\DP_OP_14_298_9081/n420 ), .Z(\DP_OP_14_298_9081/n418 ) );
  CIVXL U1817 ( .A(\DP_OP_14_298_9081/n341 ), .Z(\DP_OP_14_298_9081/n339 ) );
  CIVXL U1818 ( .A(\DP_OP_14_298_9081/n338 ), .Z(\DP_OP_14_298_9081/n337 ) );
  CIVXL U1819 ( .A(\DP_OP_14_298_9081/n448 ), .Z(\DP_OP_14_298_9081/n447 ) );
  CIVXL U1820 ( .A(\DP_OP_14_298_9081/n397 ), .Z(\DP_OP_14_298_9081/n512 ) );
  CIVXL U1821 ( .A(\DP_OP_14_298_9081/n239 ), .Z(\DP_OP_14_298_9081/n241 ) );
  CIVXL U1822 ( .A(\DP_OP_14_298_9081/n270 ), .Z(\DP_OP_14_298_9081/n268 ) );
  CIVXL U1823 ( .A(\DP_OP_14_298_9081/n457 ), .Z(\DP_OP_14_298_9081/n456 ) );
  CIVXL U1824 ( .A(\DP_OP_14_298_9081/n451 ), .Z(\DP_OP_14_298_9081/n522 ) );
  CIVXL U1825 ( .A(\DP_OP_14_298_9081/n440 ), .Z(\DP_OP_14_298_9081/n520 ) );
  COND1X1 U1826 ( .A(\DP_OP_14_298_9081/n292 ), .B(\DP_OP_14_298_9081/n1 ), 
        .C(\DP_OP_14_298_9081/n293 ), .Z(\DP_OP_14_298_9081/n2 ) );
  CND2X2 U1827 ( .A(n1496), .B(n1209), .Z(n1497) );
  COND1X2 U1828 ( .A(n1412), .B(n1629), .C(n1336), .Z(n1804) );
  COND1X1 U1829 ( .A(n1911), .B(n1809), .C(n1808), .Z(n165) );
  CENXL U1830 ( .A(n1052), .B(n1882), .Z(n1883) );
  CIVXL U1831 ( .A(n413), .Z(n1803) );
  CND2IXL U1832 ( .B(n951), .A(n1049), .Z(n1391) );
  CND2IXL U1833 ( .B(n542), .A(n1638), .Z(n1220) );
  CMXI2XL U1834 ( .A0(n1584), .A1(n1551), .S(n545), .Z(n1281) );
  CND3X1 U1835 ( .A(n1706), .B(n1731), .C(n1708), .Z(n1647) );
  CIVXL U1836 ( .A(n1731), .Z(n1733) );
  CND2XL U1837 ( .A(n1612), .B(n1422), .Z(n1613) );
  CNR2XL U1838 ( .A(n1513), .B(n1257), .Z(n1256) );
  CMXI2XL U1839 ( .A0(n1077), .A1(n1025), .S(n1411), .Z(n1850) );
  CANR1X1 U1840 ( .A(n1305), .B(n1306), .C(n1194), .Z(n1301) );
  CND2IXL U1841 ( .B(n1280), .A(n1552), .Z(n1279) );
  CNR2XL U1842 ( .A(n1669), .B(n1661), .Z(n1662) );
  CMXI2XL U1843 ( .A0(n1519), .A1(n1516), .S(n1204), .Z(n1624) );
  CNR2X2 U1844 ( .A(n1648), .B(n1647), .Z(n1702) );
  COND1XL U1845 ( .A(n1416), .B(n1925), .C(n1924), .Z(n195) );
  CANR2XL U1846 ( .A(n1923), .B(n1927), .C(n1926), .D(\C1/DATA1_1 ), .Z(n1925)
         );
  CND2XL U1847 ( .A(\C1/DATA1_0 ), .B(n1926), .Z(n1933) );
  CIVXL U1848 ( .A(n1927), .Z(n1372) );
  CANR1XL U1849 ( .A(n1356), .B(n1357), .C(n1358), .Z(n1355) );
  CND2X1 U1850 ( .A(n1183), .B(n1201), .Z(n1815) );
  CIVX2 U1851 ( .A(n1713), .Z(n1715) );
  CANR1XL U1852 ( .A(n1196), .B(\C1/DATA1_45 ), .C(n1749), .Z(n1759) );
  CNR2X1 U1853 ( .A(n1765), .B(n1761), .Z(n1750) );
  CIVX2 U1854 ( .A(n1784), .Z(n1787) );
  CND2X1 U1855 ( .A(n1183), .B(n1202), .Z(n1825) );
  CNR2X1 U1856 ( .A(n1820), .B(n1911), .Z(n1826) );
  CIVX2 U1857 ( .A(n1785), .Z(n1786) );
  CANR1XL U1858 ( .A(n1196), .B(\C1/DATA1_59 ), .C(n1682), .Z(n1690) );
  CMXI2X1 U1859 ( .A0(n1378), .A1(n1094), .S(n1425), .Z(n1765) );
  CMXI2X1 U1860 ( .A0(n1094), .A1(n1831), .S(n1425), .Z(n1842) );
  CANR1XL U1861 ( .A(n1285), .B(n1286), .C(n1422), .Z(n1284) );
  CMXI2X1 U1862 ( .A0(n1288), .A1(n1584), .S(n1206), .Z(n1287) );
  CMXI2X1 U1863 ( .A0(n1576), .A1(n1575), .S(n547), .Z(n1578) );
  CND2X1 U1864 ( .A(n1272), .B(n1193), .Z(n1271) );
  CANR1XL U1865 ( .A(n686), .B(n1612), .C(n1429), .Z(n1275) );
  CND2IX1 U1866 ( .B(n686), .A(n1265), .Z(n1264) );
  CMXI2X1 U1867 ( .A0(n1556), .A1(n1530), .S(n1206), .Z(n1265) );
  COND1XL U1868 ( .A(n542), .B(n1592), .C(n1317), .Z(n1316) );
  CANR1XL U1869 ( .A(n1318), .B(n1319), .C(n1412), .Z(n1317) );
  CIVX2 U1870 ( .A(n1720), .Z(n1381) );
  CND2X1 U1871 ( .A(n1557), .B(n1428), .Z(n1621) );
  CND2IX1 U1872 ( .B(n1426), .A(n1644), .Z(n1329) );
  CND2X1 U1873 ( .A(n1590), .B(n1425), .Z(n1854) );
  CND2IX1 U1874 ( .B(n543), .A(n1522), .Z(n1249) );
  CND2IX1 U1875 ( .B(n1485), .A(n1304), .Z(n1303) );
  CIVDX2 U1876 ( .A(n544), .Z0(n1206), .Z1(n1207) );
  CIVX3 U1877 ( .A(n544), .Z(n1424) );
  CIVX4 U1878 ( .A(n546), .Z(n1419) );
  CNIVX4 U1879 ( .A(ho_2[0]), .Z(n1418) );
  CNIVX4 U1880 ( .A(ho_2[4]), .Z(n1411) );
  CANR1XL U1881 ( .A(n1196), .B(\C1/DATA1_51 ), .C(n1386), .Z(n1382) );
  CMXI2X1 U1882 ( .A0(n1550), .A1(n1549), .S(n1419), .Z(n1584) );
  CMXI2X1 U1883 ( .A0(n1095), .A1(acc[15]), .S(n922), .Z(n1546) );
  CMXI2X1 U1884 ( .A0(acc[12]), .A1(acc[13]), .S(n922), .Z(n1539) );
  COND3XL U1885 ( .A(n1930), .B(n1929), .C(n1928), .D(n1927), .Z(n1932) );
  CENXL U1886 ( .A(n1088), .B(n1913), .Z(n1914) );
  CND2XL U1887 ( .A(n1238), .B(n1239), .Z(n1405) );
  CND2IXL U1888 ( .B(n1231), .A(n1891), .Z(n1374) );
  CENXL U1889 ( .A(n1902), .B(n1901), .Z(n1905) );
  CENXL U1890 ( .A(n1236), .B(n412), .Z(n1235) );
  CND2XL U1891 ( .A(n1217), .B(n1413), .Z(n1211) );
  CND4XL U1892 ( .A(n1786), .B(n1057), .C(n1750), .D(n1753), .Z(n1745) );
  CND2XL U1893 ( .A(n1902), .B(n1901), .Z(n1896) );
  CENXL U1894 ( .A(n1842), .B(n1841), .Z(n1845) );
  CENXL U1895 ( .A(n1737), .B(n1736), .Z(n1740) );
  CND2XL U1896 ( .A(n1057), .B(n1750), .Z(n1751) );
  CENXL U1897 ( .A(n1059), .B(n1780), .Z(n1783) );
  CENXL U1898 ( .A(n1798), .B(n1797), .Z(n1801) );
  CENXL U1899 ( .A(n1765), .B(n1764), .Z(n1768) );
  CIVXL U1900 ( .A(n1650), .Z(n1651) );
  CND2IXL U1901 ( .B(n1425), .A(n1599), .Z(n1226) );
  CMXI2XL U1902 ( .A0(acc[0]), .A1(acc[1]), .S(n922), .Z(n1322) );
  CANR1X1 U1903 ( .A(n686), .B(n1331), .C(n1194), .Z(n1330) );
  CIVXL U1904 ( .A(n1481), .Z(n1294) );
  CANR1X1 U1905 ( .A(n1280), .B(n1243), .C(n1194), .Z(n1242) );
  CIVXL U1906 ( .A(n1489), .Z(n1306) );
  CIVXL U1907 ( .A(n1493), .Z(n1608) );
  CNR2IX1 U1908 ( .B(cmd2[0]), .A(cmd2[1]), .Z(n1926) );
  CIVXL U1909 ( .A(n1334), .Z(n1930) );
  CND4XL U1910 ( .A(n1811), .B(n1413), .C(n1197), .D(n1813), .Z(n1819) );
  CIVXL U1911 ( .A(n1820), .Z(n1810) );
  COND4CX1 U1912 ( .A(n1927), .B(n1883), .C(n1199), .D(n1417), .Z(n1885) );
  CIVXL U1913 ( .A(n1057), .Z(n1762) );
  CIVXL U1914 ( .A(n1836), .Z(n1834) );
  CND3X1 U1915 ( .A(n1706), .B(n1731), .C(n1705), .Z(n1720) );
  CND2X1 U1916 ( .A(n1601), .B(n1609), .Z(n1623) );
  CND2IXL U1917 ( .B(n1206), .A(n1428), .Z(n1257) );
  CND2XL U1918 ( .A(n1206), .B(n1428), .Z(n1258) );
  CIVXL U1919 ( .A(n1557), .Z(n1331) );
  CND3X1 U1920 ( .A(n1344), .B(n1345), .C(n1346), .Z(n1520) );
  CND3X1 U1921 ( .A(n1302), .B(n1301), .C(n1303), .Z(n1510) );
  CNR2X4 U1922 ( .A(n1429), .B(n1427), .Z(n1609) );
  CEOXL U1923 ( .A(n1922), .B(n1928), .Z(n1923) );
  CIVXL U1924 ( .A(n1917), .Z(n1929) );
  CIVXL U1925 ( .A(n1796), .Z(n1744) );
  CIVXL U1926 ( .A(n1772), .Z(n1774) );
  CIVXL U1927 ( .A(n1237), .Z(n1881) );
  CNR2X1 U1928 ( .A(n1719), .B(n1911), .Z(n1718) );
  CNR2X1 U1929 ( .A(n1733), .B(n1911), .Z(n1732) );
  CNR2X1 U1930 ( .A(n1704), .B(n1911), .Z(n1703) );
  CNR2X1 U1931 ( .A(n1701), .B(n1911), .Z(n1700) );
  CND2IXL U1932 ( .B(n686), .A(n1287), .Z(n1286) );
  CMXI2X1 U1933 ( .A0(n1625), .A1(n1636), .S(n542), .Z(n1646) );
  CND2IX1 U1934 ( .B(n1203), .A(n1514), .Z(n1603) );
  CND2IX1 U1935 ( .B(n1203), .A(n1509), .Z(n1606) );
  COR2X1 U1936 ( .A(n545), .B(n686), .Z(n1348) );
  CND2IX1 U1937 ( .B(n1203), .A(n1476), .Z(n1602) );
  CND2X1 U1938 ( .A(n1486), .B(n1609), .Z(n1522) );
  CIVX4 U1939 ( .A(n1609), .Z(n1633) );
  COND4CX1 U1940 ( .A(n1933), .B(n1932), .C(n1416), .D(n1931), .Z(n196) );
  CND2X1 U1941 ( .A(n1930), .B(n1929), .Z(n1928) );
  COND4CX1 U1942 ( .A(n1367), .B(n1368), .C(n1369), .D(n1370), .Z(n186) );
  COND3X1 U1943 ( .A(n1905), .B(n1911), .C(n556), .D(n1903), .Z(n191) );
  COND4CX1 U1944 ( .A(n1337), .B(n1338), .C(n1339), .D(n1340), .Z(n184) );
  COR2X1 U1945 ( .A(n1357), .B(n1359), .Z(n1205) );
  COND4CX1 U1946 ( .A(n1880), .B(n1879), .C(n1878), .D(n1877), .Z(n183) );
  CND2X1 U1947 ( .A(n1815), .B(n1814), .Z(n1816) );
  CAOR2XL U1948 ( .A(acc[30]), .B(n1416), .C(n1195), .D(acc_a[30]), .Z(n1812)
         );
  COND3X1 U1949 ( .A(n1900), .B(n1911), .C(n555), .D(n1898), .Z(n190) );
  CAOR2XL U1950 ( .A(acc[27]), .B(n1416), .C(n1195), .D(acc_a[27]), .Z(n1843)
         );
  CAOR2XL U1951 ( .A(acc[31]), .B(n1416), .C(n1195), .D(acc_a[31]), .Z(n1807)
         );
  CAOR2XL U1952 ( .A(n918), .B(n1416), .C(n1195), .D(acc_a[47]), .Z(n1738) );
  CAOR2XL U1953 ( .A(acc[42]), .B(n1416), .C(n1195), .D(acc_a[42]), .Z(n1769)
         );
  CND2X1 U1954 ( .A(n1885), .B(n1884), .Z(n187) );
  CND2X1 U1955 ( .A(n1890), .B(n1889), .Z(n188) );
  CAOR2XL U1956 ( .A(n310), .B(n1416), .C(n1195), .D(acc_a[45]), .Z(n1749) );
  CNR2IX1 U1957 ( .B(n1707), .A(n1720), .Z(n1712) );
  CAOR2XL U1958 ( .A(acc[59]), .B(n1416), .C(n1195), .D(acc_a[59]), .Z(n1682)
         );
  CNR2X1 U1959 ( .A(n1693), .B(n1695), .Z(n1681) );
  CAOR2XL U1960 ( .A(n916), .B(n1416), .C(n1195), .D(acc_a[41]), .Z(n1781) );
  CAOR2XL U1961 ( .A(acc[16]), .B(n1416), .C(n1195), .D(acc_a[16]), .Z(n1313)
         );
  CAOR2XL U1962 ( .A(n915), .B(n1416), .C(n1195), .D(acc_a[35]), .Z(n1799) );
  CAOR2XL U1963 ( .A(n917), .B(n1416), .C(n1195), .D(acc_a[43]), .Z(n1766) );
  CND2X1 U1964 ( .A(n817), .B(n1741), .Z(n1785) );
  CNR2X1 U1965 ( .A(n1726), .B(n1911), .Z(n1728) );
  CNR2X1 U1966 ( .A(n1737), .B(n1735), .Z(n1729) );
  CNR2X1 U1967 ( .A(n1664), .B(n543), .Z(n1724) );
  CNR2X1 U1968 ( .A(n1679), .B(n1911), .Z(n1678) );
  CNR2X1 U1969 ( .A(n1833), .B(n1911), .Z(n1837) );
  CNR2X1 U1970 ( .A(n1379), .B(n306), .Z(n1248) );
  CNR2X1 U1971 ( .A(n1659), .B(n1411), .Z(n1675) );
  CND2X1 U1972 ( .A(n1743), .B(n1425), .Z(n1679) );
  CIVX2 U1973 ( .A(n1649), .Z(n1743) );
  CNR2IX1 U1974 ( .B(n1426), .A(n1742), .Z(n1685) );
  CND2X1 U1975 ( .A(n1655), .B(n1425), .Z(n1699) );
  CAOR2XL U1976 ( .A(n913), .B(n1416), .C(n1195), .D(acc_a[32]), .Z(n1362) );
  CND2X1 U1977 ( .A(n1654), .B(n1425), .Z(n1701) );
  CAN2X1 U1978 ( .A(n1644), .B(n1426), .Z(n1713) );
  CND2IX1 U1979 ( .B(n1411), .A(n1790), .Z(n1719) );
  CMXI2X1 U1980 ( .A0(n1652), .A1(n1651), .S(n543), .Z(n1653) );
  COND4CX1 U1981 ( .A(n543), .B(n1589), .C(n1284), .D(n1425), .Z(n1283) );
  CND2IX1 U1982 ( .B(n1429), .A(n1581), .Z(n1589) );
  CMXI2X1 U1983 ( .A0(n1580), .A1(n955), .S(n1427), .Z(n1581) );
  CND2X1 U1984 ( .A(n1278), .B(n1279), .Z(n1588) );
  CND2IX1 U1985 ( .B(n1429), .A(n1544), .Z(n1586) );
  CMXI2X1 U1986 ( .A0(n1543), .A1(n311), .S(n686), .Z(n1544) );
  CMXI2X1 U1987 ( .A0(n1540), .A1(n1539), .S(n1420), .Z(n1573) );
  CMXI2X1 U1988 ( .A0(n1546), .A1(n1545), .S(n1419), .Z(n1570) );
  CND2X1 U1989 ( .A(n1259), .B(n1260), .Z(n1887) );
  CND2IX1 U1990 ( .B(n1429), .A(n1533), .Z(n1591) );
  CND2IX1 U1991 ( .B(n1429), .A(n1537), .Z(n1593) );
  CMXI2X1 U1992 ( .A0(n1536), .A1(n1062), .S(n686), .Z(n1537) );
  CND2X1 U1993 ( .A(n1315), .B(n1316), .Z(n1917) );
  CMXI2X1 U1994 ( .A0(n1568), .A1(n1540), .S(n1419), .Z(n1565) );
  CND2IX1 U1995 ( .B(n1429), .A(n1564), .Z(n1592) );
  CMXI2X1 U1996 ( .A0(n1539), .A1(n1546), .S(n1420), .Z(n1560) );
  CND2IX1 U1997 ( .B(n1411), .A(n1789), .Z(n1722) );
  CIVX2 U1998 ( .A(n1735), .Z(n1705) );
  CND2IX1 U1999 ( .B(n1411), .A(n910), .Z(n1726) );
  CMXI2X1 U2000 ( .A0(n1650), .A1(n1663), .S(n543), .Z(n1742) );
  CNR2X1 U2001 ( .A(n1621), .B(n1429), .Z(n1663) );
  CND2X1 U2002 ( .A(n1622), .B(n1423), .Z(n1649) );
  CNR2X1 U2003 ( .A(n1623), .B(n543), .Z(n1660) );
  CIVX2 U2004 ( .A(n1252), .Z(n1753) );
  COAN1X1 U2005 ( .A(n1412), .B(n1620), .C(n1251), .Z(n1252) );
  CND2IX1 U2006 ( .B(n1659), .A(n541), .Z(n1251) );
  CND2X1 U2007 ( .A(n1619), .B(n1423), .Z(n1659) );
  CND2X1 U2008 ( .A(n1618), .B(n1617), .Z(n1784) );
  CND2X1 U2009 ( .A(n1412), .B(ho_2[2]), .Z(n1616) );
  CMX2X1 U2010 ( .A0(n1607), .A1(n1622), .S(n543), .Z(n1654) );
  CNR2X1 U2011 ( .A(n1606), .B(n1633), .Z(n1622) );
  CIVX2 U2012 ( .A(n1635), .Z(n1607) );
  CNR2X1 U2013 ( .A(n1603), .B(n1633), .Z(n1619) );
  COND2X1 U2014 ( .A(n1245), .B(n1244), .C(n1426), .D(n1657), .Z(n1773) );
  CMXI2X1 U2015 ( .A0(n1623), .A1(n1625), .S(n1423), .Z(n1657) );
  CNR2IX1 U2016 ( .B(n1422), .A(n1526), .Z(n1244) );
  CMXI2X1 U2017 ( .A0(n1635), .A1(n1634), .S(n1423), .Z(n1790) );
  COR2X1 U2018 ( .A(n1633), .B(n1605), .Z(n1635) );
  COR2X1 U2019 ( .A(n1633), .B(n1632), .Z(n1652) );
  CMXI2X1 U2020 ( .A0(n1627), .A1(n1637), .S(n1423), .Z(n1644) );
  COR2X1 U2021 ( .A(n1633), .B(n1604), .Z(n1627) );
  COR2X1 U2022 ( .A(n1633), .B(n1602), .Z(n1625) );
  CND2X1 U2023 ( .A(n1224), .B(n1223), .Z(n1802) );
  CMXI2X1 U2024 ( .A0(n1638), .A1(n1637), .S(n1422), .Z(n1645) );
  COR2X1 U2025 ( .A(n1633), .B(n1046), .Z(n1634) );
  COR2X1 U2026 ( .A(n1411), .B(n1599), .Z(n1327) );
  CMXI2X1 U2027 ( .A0(n1527), .A1(n946), .S(n1421), .Z(n1599) );
  CND2X1 U2028 ( .A(n1620), .B(n1411), .Z(n1326) );
  CND2X1 U2029 ( .A(n1220), .B(n1221), .Z(n1620) );
  CMXI2X1 U2030 ( .A0(n1055), .A1(n1597), .S(n1426), .Z(n1813) );
  CMXI2X1 U2031 ( .A0(n861), .A1(n1522), .S(n1422), .Z(n1830) );
  COR2X1 U2032 ( .A(n1633), .B(n1524), .Z(n1640) );
  COR2X1 U2033 ( .A(n1633), .B(n1548), .Z(n1526) );
  CND2X1 U2034 ( .A(n1600), .B(n686), .Z(n1350) );
  CND2X1 U2035 ( .A(n1519), .B(n1204), .Z(n1600) );
  CMXI2X1 U2036 ( .A0(n1515), .A1(n1527), .S(n1422), .Z(n1846) );
  CND2X1 U2037 ( .A(n1253), .B(n1254), .Z(n1527) );
  CNR2X1 U2038 ( .A(n1255), .B(n1256), .Z(n1253) );
  COR2X1 U2039 ( .A(n1633), .B(n1612), .Z(n1525) );
  CND2X1 U2040 ( .A(n1325), .B(n1324), .Z(n1222) );
  CMXI2X1 U2041 ( .A0(n1510), .A1(n1523), .S(n543), .Z(n1538) );
  CND2IX1 U2042 ( .B(n1280), .A(n1606), .Z(n1308) );
  COR2X1 U2043 ( .A(n1633), .B(n1535), .Z(n1521) );
  CMXI2X1 U2044 ( .A0(n1553), .A1(n1494), .S(n1419), .Z(n1530) );
  CND2X1 U2045 ( .A(n1230), .B(n1330), .Z(n1642) );
  CNR2X1 U2046 ( .A(n1493), .B(n1424), .Z(n1557) );
  CMXI2X1 U2047 ( .A0(n408), .A1(n1492), .S(n1203), .Z(n1229) );
  COR2X1 U2048 ( .A(n1633), .B(n1552), .Z(n1512) );
  COR2X1 U2049 ( .A(n1292), .B(n1478), .Z(n1291) );
  CND2IX1 U2050 ( .B(n686), .A(n545), .Z(n1292) );
  CND2IX1 U2051 ( .B(n1280), .A(n1604), .Z(n1290) );
  CNR2X1 U2052 ( .A(n545), .B(n686), .Z(n1293) );
  COR2X1 U2053 ( .A(n1633), .B(n1542), .Z(n1518) );
  COAN1X1 U2054 ( .A(n1348), .B(n1475), .C(n1193), .Z(n1345) );
  CND2IX1 U2055 ( .B(n1280), .A(n1602), .Z(n1344) );
  CND2X1 U2056 ( .A(n1352), .B(n1353), .Z(n1567) );
  CND2IX1 U2057 ( .B(n543), .A(n919), .Z(n1353) );
  CMXI2X1 U2058 ( .A0(n1545), .A1(n1488), .S(n1420), .Z(n1531) );
  CMXI2X1 U2059 ( .A0(acc[16]), .A1(n1069), .S(n1418), .Z(n1545) );
  CND2X1 U2060 ( .A(n920), .B(n543), .Z(n1250) );
  CMXI2X1 U2061 ( .A0(n1485), .A1(n1099), .S(n1424), .Z(n1566) );
  CND2X1 U2062 ( .A(n1242), .B(n1241), .Z(n1491) );
  CMXI2X1 U2063 ( .A0(n1445), .A1(n1439), .S(n1420), .Z(n1509) );
  CMXI2X1 U2064 ( .A0(n1442), .A1(n1438), .S(n1420), .Z(n1508) );
  CMXI2X1 U2065 ( .A0(n1474), .A1(n1437), .S(n1420), .Z(n1534) );
  CNR2IX1 U2066 ( .B(n1203), .A(n686), .Z(n1304) );
  CMXI2X1 U2067 ( .A0(n1436), .A1(n1443), .S(n1420), .Z(n1489) );
  CNR2X1 U2068 ( .A(n686), .B(n1203), .Z(n1305) );
  CMXI2X1 U2069 ( .A0(n1447), .A1(n1451), .S(n547), .Z(n1490) );
  COR2X1 U2070 ( .A(n1633), .B(n1562), .Z(n1487) );
  CMXI2X1 U2071 ( .A0(n1449), .A1(n1448), .S(n547), .Z(n1506) );
  CMXI2X1 U2072 ( .A0(n1460), .A1(n1455), .S(n547), .Z(n1503) );
  CND2IX1 U2073 ( .B(n1208), .A(n546), .Z(n1209) );
  CND2IX1 U2074 ( .B(n1465), .A(n1419), .Z(n1496) );
  COR2X1 U2075 ( .A(n1633), .B(n1559), .Z(n1641) );
  CMXI2X1 U2076 ( .A0(n1462), .A1(n1467), .S(n1419), .Z(n1502) );
  CMXI2X1 U2077 ( .A0(n1468), .A1(n1472), .S(n547), .Z(n1498) );
  CMXI2X1 U2078 ( .A0(acc[39]), .A1(acc[40]), .S(n922), .Z(n1466) );
  CMXI2X1 U2079 ( .A0(n944), .A1(n680), .S(n922), .Z(n1467) );
  CMXI2X1 U2080 ( .A0(n915), .A1(acc[36]), .S(n922), .Z(n1462) );
  CMXI2X1 U2081 ( .A0(n1465), .A1(n1464), .S(n1420), .Z(n1482) );
  CMXI2X1 U2082 ( .A0(n1069), .A1(n1063), .S(n1418), .Z(n1494) );
  CMXI2X1 U2083 ( .A0(n1514), .A1(n1511), .S(n1207), .Z(n1626) );
  CMXI2X1 U2084 ( .A0(n1459), .A1(n1208), .S(n1420), .Z(n1511) );
  CMXI2X1 U2085 ( .A0(n1458), .A1(n1457), .S(n546), .Z(n1514) );
  CMXI2X1 U2086 ( .A0(n1455), .A1(n1454), .S(n1419), .Z(n1513) );
  CIVX2 U2087 ( .A(ho_2[2]), .Z(n1423) );
  CMXI2X1 U2088 ( .A0(n1448), .A1(n1447), .S(n1420), .Z(n1517) );
  CMXI2X1 U2089 ( .A0(n1450), .A1(n1449), .S(n1420), .Z(n1473) );
  CND2IX1 U2090 ( .B(n686), .A(n1234), .Z(n1233) );
  CMXI2X1 U2091 ( .A0(n1541), .A1(n1475), .S(n1424), .Z(n1234) );
  CMXI2X1 U2092 ( .A0(n1443), .A1(n1442), .S(n1420), .Z(n1475) );
  CMXI2X1 U2093 ( .A0(acc[28]), .A1(acc[29]), .S(n1418), .Z(n1442) );
  CMXI2X1 U2094 ( .A0(n1488), .A1(n1474), .S(n1420), .Z(n1541) );
  CMXI2X1 U2095 ( .A0(n1063), .A1(acc[19]), .S(n1418), .Z(n1488) );
  CMXI2X1 U2096 ( .A0(n1437), .A1(n1436), .S(n547), .Z(n1547) );
  CMXI2X1 U2097 ( .A0(n1064), .A1(acc[23]), .S(n1418), .Z(n1437) );
  CMXI2X1 U2098 ( .A0(n1441), .A1(n1440), .S(n1420), .Z(n1516) );
  CNR2X1 U2099 ( .A(n1439), .B(n1419), .Z(n1519) );
  CMXI2X1 U2100 ( .A0(n925), .A1(acc[63]), .S(n1418), .Z(n1439) );
  CAOR2XL U2101 ( .A(n1096), .B(n1416), .C(n1195), .D(acc_a[51]), .Z(n1386) );
  CIVXL U2102 ( .A(cmd2[1]), .Z(n1433) );
  COND1XL U2103 ( .A(n1927), .B(n1876), .C(n1417), .Z(n1878) );
  CIVX2 U2104 ( .A(n542), .Z(n1421) );
  CIVXL U2105 ( .A(cmd2[0]), .Z(n1434) );
  CND3XL U2106 ( .A(n1724), .B(n1197), .C(n1425), .Z(n1665) );
  CANR1XL U2107 ( .A(n1390), .B(n1391), .C(n1392), .Z(n1389) );
  CANR1XL U2108 ( .A(n1196), .B(\C1/DATA1_24 ), .C(n1398), .Z(n1397) );
  CANR1XL U2109 ( .A(n1196), .B(\C1/DATA1_30 ), .C(n1812), .Z(n1818) );
  COND1XL U2110 ( .A(n1927), .B(n1868), .C(n1417), .Z(n1870) );
  CANR1XL U2111 ( .A(n1196), .B(\C1/DATA1_27 ), .C(n1843), .Z(n1844) );
  CANR1XL U2112 ( .A(n1196), .B(\C1/DATA1_31 ), .C(n1807), .Z(n1808) );
  CANR1XL U2113 ( .A(n1196), .B(\C1/DATA1_47 ), .C(n1738), .Z(n1739) );
  CANR1XL U2114 ( .A(n1196), .B(\C1/DATA1_42 ), .C(n1769), .Z(n1778) );
  CNR3XL U2115 ( .A(n1097), .B(n1059), .C(n937), .Z(n1770) );
  CANR1XL U2116 ( .A(n1196), .B(\C1/DATA1_41 ), .C(n1781), .Z(n1782) );
  CNR3XL U2117 ( .A(n1791), .B(n1097), .C(n937), .Z(n1779) );
  CANR1XL U2118 ( .A(n1196), .B(\C1/DATA1_16 ), .C(n1313), .Z(n1312) );
  CANR1XL U2119 ( .A(n1196), .B(\C1/DATA1_35 ), .C(n1799), .Z(n1800) );
  CANR1XL U2120 ( .A(n1196), .B(\C1/DATA1_43 ), .C(n1766), .Z(n1767) );
  CND3XL U2121 ( .A(n1727), .B(n1413), .C(n1404), .Z(n1401) );
  CAN2XL U2122 ( .A(n1726), .B(n1197), .Z(n1404) );
  COND1XL U2123 ( .A(n1911), .B(n1364), .C(n1365), .Z(n181) );
  CANR1XL U2124 ( .A(n1196), .B(\C1/DATA1_15 ), .C(n1366), .Z(n1365) );
  CANR1XL U2125 ( .A(n1196), .B(\C1/DATA1_32 ), .C(n1362), .Z(n1361) );
  CANR1XL U2126 ( .A(n686), .B(n939), .C(n1194), .Z(n1285) );
  CANR1XL U2127 ( .A(n1427), .B(n1566), .C(n1323), .Z(n1318) );
  CND3XL U2128 ( .A(n1615), .B(n1614), .C(n1613), .Z(n1618) );
  CND3XL U2129 ( .A(n1611), .B(n1423), .C(n540), .Z(n1614) );
  CANR1XL U2130 ( .A(n1411), .B(n1632), .C(n1610), .Z(n1615) );
  CND3XL U2131 ( .A(n1790), .B(n1411), .C(n1789), .Z(n1332) );
  COND1XL U2132 ( .A(n1258), .B(n948), .C(n1193), .Z(n1255) );
  CNR2IX4 U2133 ( .B(push1), .A(cmd1[1]), .Z(n202) );
  CIVX2 U2134 ( .A(n1411), .Z(n1426) );
  CIVX2 U2135 ( .A(n1411), .Z(n1425) );
  CND3XL U2136 ( .A(n1211), .B(n1213), .C(n1212), .Z(n170) );
  CND3XL U2137 ( .A(n876), .B(n1796), .C(n1752), .Z(n1755) );
  CND2XL U2138 ( .A(n1609), .B(n1616), .Z(n1610) );
  CIVXL U2139 ( .A(pushin), .Z(n1430) );
  CIVXL U2140 ( .A(pushin), .Z(n1431) );
  CIVXL U2141 ( .A(pushin), .Z(n1432) );
endmodule

